###################################################
# DK_cmos28FDSOI_6U1x_2U2x_2T8x_LB 2.1            #
###################################################
# $Id: technology.8T.12T.lef 4371 2011-10-07 11:27:22Z didier gueze $

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

UNITS
  DATABASE MICRONS 1000 ;
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  POWER MILLIWATTS 1 ;
  CURRENT MILLIAMPS 1 ;
  VOLTAGE VOLTS 1 ;
  FREQUENCY MEGAHERTZ 1 ;
END UNITS

MANUFACTURINGGRID 0.001 ;
USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
  LAYER LEF57_SPACING STRING ;
  LAYER LEF58_EOLEXTENSIONSPACING STRING ;
  LAYER LEF57_MINSTEP STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_ENCLOSUREWIDTH STRING ;
  LAYER LEF58_AREA STRING ;
  LAYER LEF58_ARRAYSPACING STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_MINIMUMCUT STRING ;
  LAYER LEF58_OPPOSITEEOLSPACING STRING ;
  LAYER LEF58_VOLTAGESPACING STRING ;
  LAYER LEF57_ANTENNAGATEPLUSDIFF STRING ;
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

##############################################################################
LAYER SLVT
##############################################################################
  TYPE IMPLANT ;
END SLVT


##############################################################################
LAYER RVT
##############################################################################
  TYPE IMPLANT ;
END RVT


##############################################################################
LAYER LVT
##############################################################################
  TYPE IMPLANT ;
END LVT


##############################################################################
LAYER DCO
##############################################################################
  TYPE IMPLANT ;
  WIDTH 0.272 ;
  SPACING 0.272 LAYER LVT ;
  SPACING 0.272 LAYER SLVT ;
  SPACING 0.272 LAYER RVT ;
END DCO

##############################################################################
LAYER NW
##############################################################################
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END NW


##############################################################################
LAYER PW
##############################################################################
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END PW


##############################################################################
LAYER PC
##############################################################################
  TYPE MASTERSLICE ;
END PC


##############################################################################
LAYER CA
##############################################################################
  TYPE    CUT ;

#  PROPERTY LEF58_ENCLOSURE "
#    ENCLOSURE ABOVE 0.006 0.006 WIDTH 0.052 EXCEPTEXTRACUT 0.060 ;
#    ENCLOSURE ABOVE 0.000 0.000 WIDTH 0.053 ;
#  " ; # 505b

END CA


##############################################################################
LAYER M1
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   VERTICAL ;
  PITCH       0.136 0.100 ;
  OFFSET      0.068 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 500
  MAXWIDTH    4.500 ; # 500b

  #SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes
  SPACING 0.069 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 502, 504

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES R 504k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
      ENDOFLINE 0.058 EXTENSION 0.01
      ENDOFLINE 0.105 EXTENSION 0.008 ENDTOEND 0.006
      MINLENGTH 0.041 TWOSIDES ;
  " ; # ALP5_502

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.041
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    EXCEPTEDGELENGTH 0.072 PRL 0.01
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 506a 506b 506c 506d

  AREA                  0.0093 ; # 501a
  PROPERTY LEF58_AREA "
    AREA 0.010 EXCEPTMINSIZE 0.072 0.072 ;
    AREA 0.030 EXCEPTEDGELENGTH 0.13 ;
  " ; # 501aSE  501d
  MINENCLOSEDAREA       0.048 ; # 501b

  MINSTEP 0.049 MAXEDGES 1 ; # SE4

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 FROMABOVE ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 FROMABOVE ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE AREA 0.0338 WITHIN 1.001 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.000 FROMABOVE AREA 0.9999 WITHIN 2.101 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.800 FROMABOVE AREA 8.9999 WITHIN 5.501 ;
  " ; # 612abc 613abc

## 502j1, 502j2, 502j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M1


##############################################################################
LAYER V1
##############################################################################

  TYPE    CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS VX    WIDTH 0.050 ;
    CUTCLASS VXBAR WIDTH 0.050 LENGTH 0.100 CUTS 2 ;
    CUTCLASS VXLRG WIDTH 0.100 LENGTH 0.100 CUTS 2 ;
  " ; # 550 550b 550c 550d 612b2

  PROPERTY LEF58_ENCLOSUREWIDTH "
    ENCLOSUREWIDTH VIAOVERLAPONLY ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS VX 0.008 0.008 ;
    ENCLOSURE CUTCLASS VX BELOW 0.011 0.003 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VX BELOW 0.011 0.003 WIDTH 0.050 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 WIDTH 0.082 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.082 ;
    ENCLOSURE CUTCLASS VX BELOW 0.011 0.003 WIDTH 0.082 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX BELOW 0.000 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.005 0.005 WIDTH 0.085 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.010 0.010 WIDTH 0.100 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.014 WIDTH 0.143 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VXLRG 0.017 0.017 ;
    ENCLOSURE CUTCLASS VXBAR END 0.017 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.008 SIDE 0.008 WIDTH 0.073 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.010 SIDE 0.010 WIDTH 0.105 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.014 SIDE 0.014 WIDTH 0.143 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.026 SIDE 0.025 WIDTH 0.151 ;
  " ; # 570a,b,c 571a,b,c 572_or 572a,b,c,d 610 611 615 615c 675c

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             0.134 0.134   0.080 0.080   0.080 0.080   0.100 0.100
      VXLRG          0.080 0.080   0.100 0.100   0.080 0.080   0.080 0.080
      VXBAR SIDE     0.080 0.080   0.080 0.080   0.076 0.076   0.103 0.103
      VXBAR END      0.100 0.100   0.080 0.080   0.103 0.103   0.130 0.130 ;
  " ; # 553 553bb 553c 553d 553e 553f 553g 553h 553i 553q

  PROPERTY LEF58_SPACING "
    SPACING 0.141 CENTERTOCENTER ADJACENTCUTS 2 EXACTALIGNED 3 WITHIN 0.141 CUTCLASS VX ;
  " ; # 553q1,q2

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END V1


##############################################################################
LAYER M2
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       0.100 0.100 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 600
  MAXWIDTH    4.500 ; # 600b

  SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 602, 604

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES 604k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
    ENDOFLINE 0.105 EXTENSION 0.010
    MINLENGTH 0.021 TWOSIDES ; " ; # ALP5_602a

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.021
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 606a 606b 606c 606d

  AREA                  0.011 ; # 601a
  PROPERTY LEF58_AREA "AREA 0.030 EXCEPTEDGELENGTH 0.13 ;" ; # 601aSE
  MINENCLOSEDAREA       0.059 ; # 601b

  MINSTEP 0.050 MAXEDGES 1 ; # SE5

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 WITHIN 2 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW LENGTH 0.184 WITHIN 0.005 ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE AREA 0.0338 WITHIN 1.001 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.000 FROMABOVE AREA 0.9999 WITHIN 2.101 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.800 FROMABOVE AREA 8.9999 WITHIN 5.501 ;
  " ; # 612abc 613abc

## 602i1, 602i2, 602i4 602j1, 602j2, 602j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M2


##############################################################################
LAYER V2
##############################################################################

  TYPE    CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS VX    WIDTH 0.050 ;
    CUTCLASS VXBAR WIDTH 0.050 LENGTH 0.100 CUTS 2 ;
    CUTCLASS VXLRG WIDTH 0.100 LENGTH 0.100 CUTS 2 ;
  " ; # 550 550b 550c 550d

  PROPERTY LEF58_ENCLOSUREWIDTH "
    ENCLOSUREWIDTH VIAOVERLAPONLY ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS VX 0.008 0.008 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX 0.008 0.008 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.073 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.010 0.010 WIDTH 0.105 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.014 WIDTH 0.143 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VXLRG 0.017 0.017 ;
    ENCLOSURE CUTCLASS VXBAR END 0.017 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.008 SIDE 0.008 WIDTH 0.073 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.010 SIDE 0.010 WIDTH 0.105 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.014 SIDE 0.014 WIDTH 0.143 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.026 SIDE 0.025 WIDTH 0.151 ;
  " ; # 570a,b,c 571a,b,c 572_or 572a,b,c,d 610 611 615 615c 675c

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             0.134 0.134   0.080 0.080   0.080 0.080   0.100 0.100
      VXLRG          0.080 0.080   0.100 0.100   0.080 0.080   0.080 0.080
      VXBAR SIDE     0.080 0.080   0.080 0.080   0.076 0.076   0.103 0.103
      VXBAR END      0.100 0.100   0.080 0.080   0.103 0.103   0.130 0.130 ;
  " ; # 553 553bb 553c 553d 553e 553f 553g 553h 553i 553q

  PROPERTY LEF58_SPACING "
    SPACING 0.141 CENTERTOCENTER ADJACENTCUTS 2 EXACTALIGNED 3 WITHIN 0.141 CUTCLASS VX ;
  " ; # 553q1,q2

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      LAYER V1
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX           0.115 0.115     0.144 0.144   0.069 0.069   0.069 0.069
      VXLRG        0.144 0.144     0 0           0.069 0.069   0.069 0.069
      VXBAR SIDE   0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069
      VXBAR END    0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069 ;
    SPACINGTABLE
      DEFAULT 0
      SAMENET
      LAYER V1
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             - -           - -           - -           - -
      VXLRG          - -           - -           - -           - -
      VXBAR SIDE     - -           - -           - -           - -
      VXBAR END      - -           - -           - -           - - ;
  " ; # 555b 555d 555dd 555e 555i

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END V2


##############################################################################
LAYER M3
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   VERTICAL ;
  PITCH       0.100 0.100 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 600
  MAXWIDTH    4.500 ; # 600b

  SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 602, 604

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES 604k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
    ENDOFLINE 0.105 EXTENSION 0.010
    MINLENGTH 0.021 TWOSIDES ;
  " ; # ALP5_602a

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.021
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 606a 606b 606c 606d

  AREA                  0.011 ; # 601a
  PROPERTY LEF58_AREA "AREA 0.030 EXCEPTEDGELENGTH 0.13 ;" ; # 601aSE
  MINENCLOSEDAREA       0.059 ; # 601b

  MINSTEP 0.050 MAXEDGES 1 ; # SE5

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW LENGTH 0.184 WITHIN 0.005 ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE AREA 0.0338 WITHIN 1.001 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.000 FROMABOVE AREA 0.9999 WITHIN 2.101 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.800 FROMABOVE AREA 8.9999 WITHIN 5.501 ;
  " ; # 612abc 613abc

## 602i1, 602i2, 602i4 602j1, 602j2, 602j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M3


##############################################################################
LAYER V3
##############################################################################

  TYPE    CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS VX    WIDTH 0.050 ;
    CUTCLASS VXBAR WIDTH 0.050 LENGTH 0.100 CUTS 2 ;
    CUTCLASS VXLRG WIDTH 0.100 LENGTH 0.100 CUTS 2 ;
  " ; # 550 550b 550c 550d

  PROPERTY LEF58_ENCLOSUREWIDTH "
    ENCLOSUREWIDTH VIAOVERLAPONLY ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS VX 0.008 0.008 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX 0.008 0.008 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.073 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.010 0.010 WIDTH 0.105 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.014 WIDTH 0.143 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VXLRG 0.017 0.017 ;
    ENCLOSURE CUTCLASS VXBAR END 0.017 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.008 SIDE 0.008 WIDTH 0.073 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.010 SIDE 0.010 WIDTH 0.105 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.014 SIDE 0.014 WIDTH 0.143 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.026 SIDE 0.025 WIDTH 0.151 ;
  " ; # 570a,b,c 571a,b,c 572_or 572a,b,c,d 610 611 615 615c 675c

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             0.134 0.134   0.080 0.080   0.080 0.080   0.100 0.100
      VXLRG          0.080 0.080   0.100 0.100   0.080 0.080   0.080 0.080
      VXBAR SIDE     0.080 0.080   0.080 0.080   0.076 0.076   0.103 0.103
      VXBAR END      0.100 0.100   0.080 0.080   0.103 0.103   0.130 0.130 ;
  " ; # 553 553bb 553c 553d 553e 553f 553g 553h 553i 553q

  PROPERTY LEF58_SPACING "
    SPACING 0.141 CENTERTOCENTER ADJACENTCUTS 2 EXACTALIGNED 3 WITHIN 0.141 CUTCLASS VX ;
  " ; # 553q1,q2

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      LAYER V2
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX           0.115 0.115     0.144 0.144   0.069 0.069   0.069 0.069
      VXLRG        0.144 0.144     0 0           0.069 0.069   0.069 0.069
      VXBAR SIDE   0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069
      VXBAR END    0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069 ;
    SPACINGTABLE
      DEFAULT 0
      SAMENET
      LAYER V2
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             - -           - -           - -           - -
      VXLRG          - -           - -           - -           - -
      VXBAR SIDE     - -           - -           - -           - -
      VXBAR END      - -           - -           - -           - - ;
  " ; # 555b 555d 555dd 555e 555i

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END V3


##############################################################################
LAYER M4
##############################################################################
  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       0.100 0.100 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 600
  MAXWIDTH    4.500 ; # 600b

  SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 602, 604

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES 604k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
    ENDOFLINE 0.105 EXTENSION 0.010
    MINLENGTH 0.021 TWOSIDES ; " ; # ALP5_602a

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.021
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 606a 606b 606c 606d

  AREA                  0.011 ; # 601a
  PROPERTY LEF58_AREA "AREA 0.030 EXCEPTEDGELENGTH 0.13 ;" ; # 601aSE
  MINENCLOSEDAREA       0.059 ; # 601b

  MINSTEP 0.050 MAXEDGES 1 ; # SE5

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW LENGTH 0.184 WITHIN 0.005 ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE AREA 0.0338 WITHIN 1.001 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.000 FROMABOVE AREA 0.9999 WITHIN 2.101 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.800 FROMABOVE AREA 8.9999 WITHIN 5.501 ;
  " ; # 612abc 613abc

## 602i1, 602i2, 602i4 602j1, 602j2, 602j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M4


##############################################################################
LAYER V4
##############################################################################

  TYPE    CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS VX    WIDTH 0.050 ;
    CUTCLASS VXBAR WIDTH 0.050 LENGTH 0.100 CUTS 2 ;
    CUTCLASS VXLRG WIDTH 0.100 LENGTH 0.100 CUTS 2 ;
  " ; # 550 550b 550c 550d

  PROPERTY LEF58_ENCLOSUREWIDTH "
    ENCLOSUREWIDTH VIAOVERLAPONLY ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS VX 0.008 0.008 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX 0.008 0.008 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.073 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.010 0.010 WIDTH 0.105 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.014 WIDTH 0.143 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VXLRG 0.017 0.017 ;
    ENCLOSURE CUTCLASS VXBAR END 0.017 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.008 SIDE 0.008 WIDTH 0.073 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.010 SIDE 0.010 WIDTH 0.105 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.014 SIDE 0.014 WIDTH 0.143 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.026 SIDE 0.025 WIDTH 0.151 ;
  " ; # 570a,b,c 571a,b,c 572_or 572a,b,c,d 610 611 615 615c 675c

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             0.134 0.134   0.080 0.080   0.080 0.080   0.100 0.100
      VXLRG          0.080 0.080   0.100 0.100   0.080 0.080   0.080 0.080
      VXBAR SIDE     0.080 0.080   0.080 0.080   0.076 0.076   0.103 0.103
      VXBAR END      0.100 0.100   0.080 0.080   0.103 0.103   0.130 0.130 ;
  " ; # 553 553bb 553c 553d 553e 553f 553g 553h 553i 553q

  PROPERTY LEF58_SPACING "
    SPACING 0.141 CENTERTOCENTER ADJACENTCUTS 2 EXACTALIGNED 3 WITHIN 0.141 CUTCLASS VX ;
  " ; # 553q1,q2

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      LAYER V3
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX           0.115 0.115     0.144 0.144   0.069 0.069   0.069 0.069
      VXLRG        0.144 0.144     0 0           0.069 0.069   0.069 0.069
      VXBAR SIDE   0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069
      VXBAR END    0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069 ;
    SPACINGTABLE
      DEFAULT 0
      SAMENET
      LAYER V3
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             - -           - -           - -           - -
      VXLRG          - -           - -           - -           - -
      VXBAR SIDE     - -           - -           - -           - -
      VXBAR END      - -           - -           - -           - - ;
  " ; # 555b 555d 555dd 555e 555i

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END V4


##############################################################################
LAYER M5
##############################################################################
  TYPE        ROUTING ;
  DIRECTION   VERTICAL ;
  PITCH       0.100 0.100 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 600
  MAXWIDTH    4.500 ; # 600b

  SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 602, 604

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES 604k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
    ENDOFLINE 0.105 EXTENSION 0.010
    MINLENGTH 0.021 TWOSIDES ; " ; # ALP5_602a

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.021
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 606a 606b 606c 606d

  AREA                  0.011 ; # 601a
  PROPERTY LEF58_AREA "AREA 0.030 EXCEPTEDGELENGTH 0.13 ;" ; # 601aSE
  MINENCLOSEDAREA       0.059 ; # 601b

  MINSTEP 0.050 MAXEDGES 1 ; # SE5

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW LENGTH 0.184 WITHIN 0.005 ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMABOVE AREA 0.0338 WITHIN 1.001 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.000 FROMABOVE AREA 0.9999 WITHIN 2.101 ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 1.800 FROMABOVE AREA 8.9999 WITHIN 5.501 ;
  " ; # 612abc 613abc

## 602i1, 602i2, 602i4 602j1, 602j2, 602j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M5


##############################################################################
LAYER V5
##############################################################################

  TYPE    CUT ;

  PROPERTY LEF58_CUTCLASS "
    CUTCLASS VX    WIDTH 0.050 ;
    CUTCLASS VXBAR WIDTH 0.050 LENGTH 0.100 CUTS 2 ;
    CUTCLASS VXLRG WIDTH 0.100 LENGTH 0.100 CUTS 2 ;
  " ; # 550 550b 550c 550d

  PROPERTY LEF58_ENCLOSUREWIDTH "
    ENCLOSUREWIDTH VIAOVERLAPONLY ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS VX 0.008 0.008 ;
    ENCLOSURE CUTCLASS VX BELOW 0.017 0.000 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 EXTRACUT ;
    ENCLOSURE CUTCLASS VX 0.008 0.008 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX ABOVE 0.032 0.000 REDUNDANTCUT 0.226 ;
    ENCLOSURE CUTCLASS VX BELOW 0.008 0.008 WIDTH 0.073 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.010 0.010 WIDTH 0.105 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VX BELOW 0.014 0.014 WIDTH 0.143 EXCEPTEXTRACUT 0.226 PRL ;
    ENCLOSURE CUTCLASS VXLRG 0.017 0.017 ;
    ENCLOSURE CUTCLASS VXBAR END 0.017 SIDE 0.000 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.008 SIDE 0.008 WIDTH 0.073 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.010 SIDE 0.010 WIDTH 0.105 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.014 SIDE 0.014 WIDTH 0.143 ;
    ENCLOSURE CUTCLASS VXBAR BELOW END 0.026 SIDE 0.025 WIDTH 0.151 ;
  " ; # 570a,b,c 571a,b,c 572_or 572a,b,c,d 610 611 615 615c 675c

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             0.134 0.134   0.080 0.080   0.080 0.080   0.100 0.100
      VXLRG          0.080 0.080   0.100 0.100   0.080 0.080   0.080 0.080
      VXBAR SIDE     0.080 0.080   0.080 0.080   0.076 0.076   0.103 0.103
      VXBAR END      0.100 0.100   0.080 0.080   0.103 0.103   0.130 0.130 ;
  " ; # 553 553bb 553c 553d 553e 553f 553g 553h 553i 553q

  PROPERTY LEF58_SPACING "
    SPACING 0.141 CENTERTOCENTER ADJACENTCUTS 2 EXACTALIGNED 3 WITHIN 0.141 CUTCLASS VX ;
  " ; # 553q1,q2

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      LAYER V4
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX           0.115 0.115     0.144 0.144   0.069 0.069   0.069 0.069
      VXLRG        0.144 0.144     0 0           0.069 0.069   0.069 0.069
      VXBAR SIDE   0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069
      VXBAR END    0.069 0.069     0.069 0.069   0.069 0.069   0.069 0.069 ;
    SPACINGTABLE
      DEFAULT 0
      SAMENET
      LAYER V4
      CENTERTOCENTER VX TO VX
      CUTCLASS       VX            VXLRG         VXBAR SIDE    VXBAR END
      VX             - -           - -           - -           - -
      VXLRG          - -           - -           - -           - -
      VXBAR SIDE     - -           - -           - -           - -
      VXBAR END      - -           - -           - -           - - ;
  " ; # 555b 555d 555dd 555e 555i

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END V5


##############################################################################
LAYER M6
##############################################################################
  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       0.100 0.100 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.050 ;
  MINWIDTH    0.050 ; # 600
  MAXWIDTH    4.500 ; # 600b

  SPACING 0.100 NOTCHLENGTH 0.075 ; # Avoid U-shapes

  SPACINGTABLE  TWOWIDTHS
                 # WIDTH    0.000  0.072  0.156  0.208  0.700  1.500
                 # PRL      0.000  0.000  0.000  0.300  0.700  1.500
                 # -------------------------------------------------
    WIDTH 0.000             0.050  0.050  0.066  0.095  0.165  0.500
    WIDTH 0.072  PRL 0.000  0.050  0.050  0.074  0.103  0.173  0.500
    WIDTH 0.156  PRL 0.000  0.066  0.074  0.082  0.111  0.181  0.500
    WIDTH 0.208  PRL 0.300  0.095  0.103  0.111  0.140  0.210  0.500
    WIDTH 0.700  PRL 0.700  0.165  0.173  0.181  0.210  0.280  0.500
    WIDTH 1.500  PRL 1.500  0.500  0.500  0.500  0.500  0.500  0.500 ; # 602, 604

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      PARALLELSPANLENGTH  PRL 0.104
      SPANLENGTH      0       0.05    0.058   0.059   0.062
      SPANLENGTH      0.072   0.058   0.065   0.065   0.065
      SPANLENGTH      0.156   0.059   0.065   0.068   0.068
      SPANLENGTH      0.208   0.062   0.065   0.068   0.074 ;
  " ; # SPAN RULES 604k-m

  PROPERTY LEF58_EOLEXTENSIONSPACING "
    EOLEXTENSIONSPACING 0.05
    ENDOFLINE 0.105 EXTENSION 0.010
    MINLENGTH 0.021 TWOSIDES ; " ; # ALP5_602a

  PROPERTY LEF58_OPPOSITEEOLSPACING "
    OPPOSITEEOLSPACING
    WIDTH 0.065
    ENDWIDTH 0.105 MINLENGTH 0.021
    JOINTLENGTH 0.072 JOINTTOEDGEEND 0.070
    ENDTOEND 0.065 0.070
    ENDTOJOINT 0.065 0.065
    JOINTTOEND 0.060 0.070
    JOINTTOJOINT 0.060 0.070 ;
  " ; # 606a 606b 606c 606d

  AREA                  0.011 ; # 601a
  PROPERTY LEF58_AREA "AREA 0.030 EXCEPTEDGELENGTH 0.13 ;" ; # 601aSE
  MINENCLOSEDAREA       0.059 ; # 601b

  MINSTEP 0.050 MAXEDGES 1 ; # SE5

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW ;
    MINIMUMCUT CUTCLASS VX 2 WIDTH 0.184 FROMBELOW LENGTH 0.184 WITHIN 0.005 ;
    MINIMUMCUT CUTCLASS VX 3 CUTCLASS VXLRG 2 CUTCLASS VXBAR 2 WIDTH 0.330 FROMBELOW ;
    MINIMUMCUT CUTCLASS VX 4 CUTCLASS VXLRG 3 CUTCLASS VXBAR 3 WIDTH 0.460 FROMBELOW ;
  " ; # 612abc 613abc

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT 2 WIDTH 0.345 FROMABOVE ;
    MINIMUMCUT 3 WIDTH 0.545 FROMABOVE ;
    MINIMUMCUT 4 WIDTH 0.745 FROMABOVE ;
    MINIMUMCUT 2 WIDTH 0.700 FROMABOVE AREA  0.4899 WITHIN 1.401 ;
    MINIMUMCUT 2 WIDTH 2.000 FROMABOVE AREA  3.9999 WITHIN 2.801 ;
    MINIMUMCUT 2 WIDTH 3.000 FROMABOVE AREA 29.9999 WITHIN 7.101 ;
  " ; # 2x72a, 2x72ab, 2x72b, 2x72bb, 2x72c, 2x72cb, 2x73a, 2x73b, 2x73c

## 602i1, 602i2, 602i4 602j1, 602j2, 602j4
# PROPERTY LEF58_VOLTAGESPACING "
#   VOLTAGESPACING TOCUT ABOVE
#      1.5   0.070
#      1.8   0.090
#      2.5   0.125
#      3.3   0.165 ;
# " ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END M6


##############################################################################
LAYER W0
##############################################################################

  TYPE    CUT ;

  WIDTH   0.100 ; # 2x50
  SPACING 0.230 CENTERTOCENTER ; # 2x53b
  SPACING 0.250 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.250 ; # 2x53a
  SPACING 0.100 SAMENET ; # 2x53

  PROPERTY LEF58_ARRAYSPACING "
    ARRAYSPACING PARALLELOVERLAP LONGARRAY CUTSPACING 0.100
      ARRAYCUTS 4 SPACING 0.300
      ARRAYCUTS 5 SPACING 0.500
      ARRAYCUTS 6 SPACING 0.700 ;
  " ; # 2x51a, 2x51b, 2x51c, 2x51d

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE LAYER V5 CENTERTOCENTER ALL TO VX
    CUTCLASS         ALL
    VX           0.155 0.155
    VXLRG        0.182 0.182
    VXBAR SIDE   0.082 0.082
    VXBAR END    0.082 0.082 ;
      SPACINGTABLE
       DEFAULT 0
       SAMENET
       LAYER V5
       CENTERTOCENTER ALL TO VX
       CUTCLASS       ALL
       VX             - -
       VXLRG          - -
       VXBAR SIDE     - -
       VXBAR END      - - ;
  " ; # 555j,k,l

  ENCLOSURE BELOW 0.020 0.020 ; # 2x60a
  ENCLOSURE BELOW 0.030 0.010 ; # 2x60b
  ENCLOSURE BELOW 0.040 0.000 ; # 2x60c
  ENCLOSURE ABOVE 0.020 0.020 ; # 2x61a
  ENCLOSURE ABOVE 0.030 0.010 ; # 2x61b
  ENCLOSURE ABOVE 0.040 0.000 ; # 2x61c
  ENCLOSURE BELOW 0.015 0.015 WIDTH 0.179 EXCEPTEXTRACUT 0.129 ; # 2x60f
  ENCLOSURE BELOW 0.035 0.035 WIDTH 0.490 ; # 2x73 Note nr 2 !!!

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END W0


##############################################################################
LAYER B1
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   VERTICAL ;
  PITCH       0.200 0.200 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.100 ;
  MINWIDTH    0.100 ; # 2x00
  MAXWIDTH    12.000 ; # 2x00b

  SPACINGTABLE  TWOWIDTHS
                     # WIDTH    0.000  0.315  1.000  1.500  4.500
                     # PRL      0.000  0.000  0.000  1.500  4.500
                     # ------------------------------------------
    WIDTH 0.000                 0.100  0.145  0.250  0.250  0.250
    WIDTH 0.315    PRL 0.000    0.145  0.200  0.300  0.300  0.300
    WIDTH 1.000    PRL 0.000    0.250  0.300  0.400  0.400  0.400
    WIDTH 1.500    PRL 1.500    0.250  0.300  0.400  0.500  0.500
    WIDTH 4.500    PRL 4.500    0.250  0.300  0.400  0.500  1.500 ; # 2x02, 2x04, 2x04a, 2x04b, 2x04c, 2x04d, 2x04e, 2x04f

  AREA                  0.040 ; # 2x01a
  MINENCLOSEDAREA       0.135 ; # 2x01b

  MINSTEP 0.100 MAXEDGES 1 ; # SE7

  MINIMUMCUT 2 WIDTH 0.345 ; # 2x72a, 2x72ab
  MINIMUMCUT 3 WIDTH 0.545 ; # 2x72b, 2x72bb
  MINIMUMCUT 4 WIDTH 0.745 ; # 2x72c, 2x72cb

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT 2 WIDTH 0.700 AREA  0.4899 WITHIN 1.401 ;
    MINIMUMCUT 2 WIDTH 2.000 AREA  3.9999 WITHIN 2.801 ;
    MINIMUMCUT 2 WIDTH 3.000 AREA 29.9999 WITHIN 7.101 ;
  " ; # 2x73a, 2x73b, 2x73c

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END B1


##############################################################################
LAYER W1
##############################################################################

  TYPE    CUT ;

  WIDTH   0.100 ; # 2x50
  SPACING 0.230 CENTERTOCENTER ; # 2x53b
  SPACING 0.250 CENTERTOCENTER ADJACENTCUTS 3 WITHIN 0.250 ; # 2x53a
  SPACING 0.100 SAMENET ; # 2x53

  PROPERTY LEF58_ARRAYSPACING "
    ARRAYSPACING PARALLELOVERLAP LONGARRAY CUTSPACING 0.100
      ARRAYCUTS 4 SPACING 0.300
      ARRAYCUTS 5 SPACING 0.500
      ARRAYCUTS 6 SPACING 0.700 ;
  " ; # 2x51a, 2x51b, 2x51c, 2x51d

  ENCLOSURE BELOW 0.020 0.020 ; # 2x62a
  ENCLOSURE BELOW 0.030 0.010 ; # 2x62b
  ENCLOSURE BELOW 0.040 0.000 ; # 2x62c
  ENCLOSURE ABOVE 0.020 0.020 ; # 2x63a
  ENCLOSURE ABOVE 0.030 0.010 ; # 2x63b
  ENCLOSURE ABOVE 0.040 0.000 ; # 2x63c
  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE BELOW 0.015 0.015 WIDTH 0.180 EXCEPTEXTRACUT 0.300 ;
    ENCLOSURE BELOW 0.020 0.020 WIDTH 0.296 EXCEPTEXTRACUT 0.300 PRL ;
    ENCLOSURE BELOW 0.068 0.068 WIDTH 0.776 EXCEPTEXTRACUT 0.300 PRL ;
  " ; # 2x62f 2x75a 2x75b


  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END W1


##############################################################################
LAYER B2
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       0.200 0.200 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.100 ;
  MINWIDTH    0.100 ; # 2x00
  MAXWIDTH    12.000 ; # 2x00b

  SPACINGTABLE  TWOWIDTHS
                     # WIDTH    0.000  0.315  1.000  1.500  4.500
                     # PRL      0.000  0.000  0.000  1.500  4.500
                     # ------------------------------------------
    WIDTH 0.000                 0.100  0.145  0.250  0.250  0.250
    WIDTH 0.315    PRL 0.000    0.145  0.200  0.300  0.300  0.300
    WIDTH 1.000    PRL 0.000    0.250  0.300  0.400  0.400  0.400
    WIDTH 1.500    PRL 1.500    0.250  0.300  0.400  0.500  0.500
    WIDTH 4.500    PRL 4.500    0.250  0.300  0.400  0.500  1.500 ; # 2x02, 2x04, 2x04a, 2x04b, 2x04c, 2x04d, 2x04e, 2x04f

  AREA                  0.040 ; # 2x01a
  MINENCLOSEDAREA       0.135 ; # 2x01b

  MINSTEP 0.100 MAXEDGES 1 ; # SE7

  MINIMUMCUT 2 WIDTH 0.345 FROMBELOW ; # 2x72a, 2x72ab
  MINIMUMCUT 3 WIDTH 0.545 FROMBELOW ; # 2x72b, 2x72bb
  MINIMUMCUT 4 WIDTH 0.745 FROMBELOW ; # 2x72c, 2x72cb

  PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT 2 WIDTH 0.700 FROMBELOW AREA  0.4899 WITHIN 1.401 ;
    MINIMUMCUT 2 WIDTH 2.000 FROMBELOW AREA  3.9999 WITHIN 2.801 ;
    MINIMUMCUT 2 WIDTH 3.000 FROMBELOW AREA 29.9999 WITHIN 7.101 ;
  " ; # 2x73a, 2x73b, 2x73c

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END B2


##############################################################################
LAYER YZ
##############################################################################

  TYPE    CUT ;

  WIDTH   0.360 ; # 8x50_YZ
  SPACING 0.440 ; # 8x53_YZ

  ENCLOSURE BELOW 0.080 0.020 ; # 8x60a_YZ, 8x60_YZ
  ENCLOSURE ABOVE 0.080 0.020 ; # 8x61_YZ, 8x61a_YZ

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END YZ


##############################################################################
LAYER IA
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       0.800 0.800 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.400 ;
  MINWIDTH    0.400 ; # 8x00
  MAXWIDTH    12.000 ; # 8x00b

  SPACINGTABLE  TWOWIDTHS
                   # WIDTH    0.000  2.000  4.000  8.000
                   # PRL      0.000  2.000  4.000  8.000
                   # -----------------------------------
  WIDTH 0.000                 0.400  0.600  1.000  2.000
  WIDTH 2.000    PRL 2.000    0.600  0.800  1.200  2.000
  WIDTH 4.000    PRL 4.000    1.000  1.200  1.600  2.000
  WIDTH 8.000    PRL 8.000    2.000  2.000  2.000  4.000 ; # 8x04, 8x04a, 8x04b, 8x04c, 8x04d, 8x04e, 8x04f

  AREA                  0.480 ; # 8x01a
  MINENCLOSEDAREA       0.870 ; # 8x01b

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END IA


##############################################################################
LAYER XA
##############################################################################

  TYPE    CUT ;

  WIDTH   0.360 ; # 8Bx50
  SPACING 0.440 SAMENET ; # R 8Bx53
  SPACING 0.560 ; # R 8Bx53b

  ENCLOSURE BELOW 0.080 0.020 ; # 8Bx62, 8Bx62a
  ENCLOSURE ABOVE 0.080 0.020 ; # 8Bx63, 8Bx63a

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 5.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END XA


##############################################################################
LAYER IB
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   VERTICAL ;
  PITCH       0.800 0.800 ;
  OFFSET      0.000 0.000 ;
  WIDTH       0.400 ;
  MINWIDTH    0.400 ; # 8x00
  MAXWIDTH    12.000 ; # 8x00b

  SPACINGTABLE  TWOWIDTHS
                   # WIDTH    0.000  2.000  4.000  8.000
                   # PRL      0.000  2.000  4.000  8.000
                   # -----------------------------------
  WIDTH 0.000                 0.400  0.600  1.000  2.000
  WIDTH 2.000    PRL 2.000    0.600  0.800  1.200  2.000
  WIDTH 4.000    PRL 4.000    1.000  1.200  1.600  2.000
  WIDTH 8.000    PRL 8.000    2.000  2.000  2.000  4.000 ; # 8x04, 8x04a, 8x04b, 8x04c, 8x04d, 8x04e, 8x04f

  AREA                  0.480 ; # 8x01a
  MINENCLOSEDAREA       0.870 ; # 8x01b

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 2000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 500.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;
  ANTENNAMODEL OXIDE3 ;
  ANTENNADIFFAREARATIO 150.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 50.0 ;" ;

END IB


##############################################################################
LAYER VV
##############################################################################

  TYPE    CUT ;

  WIDTH   3.000 ; # LB50
  SPACING 2.000 ; # LB53

  ENCLOSURE BELOW 0.500 0.500 ; # LB70
  ENCLOSURE ABOVE 1.000 1.000 ; # LB75

END VV


##############################################################################
LAYER LB
##############################################################################

  TYPE        ROUTING ;
  DIRECTION   HORIZONTAL ;
  PITCH       10.000 10.000 ;
  OFFSET      0.000 0.000 ;
  WIDTH       4.000 ;
  MINWIDTH    4.000 ; # LB00
  MAXWIDTH    35.000 ; # LB.W.2
  SPACING     2.000 ; # LB02

# The rule LB04b only applies in flip chip and not in wiremode
# Wiremode is currently not supported in the DPs
#  SPACINGTABLE  TWOWIDTHS
#                 # WIDTH    0.000  35.000
#                 # ----------------------
#    WIDTH  0.000            2.000   4.000
#    WIDTH 35.000            4.000   4.000 ; # LB02, LB04b

END LB


##############################################################################
LAYER overlap
##############################################################################
  TYPE OVERLAP ;
END overlap


################################## VIA FOR ROUTING ######################################
# Automatically generated by generateViaLEF

VIA CDS_V12_1x1_SV DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.033  0.033  0.033 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V12_1x1_SV

VIA CDS_V12_1x1_SH DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.033  0.033  0.033 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V12_1x1_SH

VIA CDS_V12_1x1_VH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V12_1x1_VH

VIA CDS_V12_1x1_VV DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V12_1x1_VV

VIA CDS_V12_1x1_HH DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V12_1x1_HH

VIA CDS_V12_1x1_HV DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V12_1x1_HV

VIA CDS_V12_1x2_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V1 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M2 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V12_1x2_CENTER

VIA CDS_V12_1x2_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V12_1x2_NORTH

VIA CDS_V12_1x2_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V1 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V12_1x2_SOUTH

VIA CDS_V12_2x1_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.092 -0.039  0.092  0.039 ;
  LAYER V1 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M2 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V12_2x1_CENTER

VIA CDS_V12_2x1_EAST DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.039  0.159  0.039 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V12_2x1_EAST

VIA CDS_V12_2x1_WEST DEFAULT
  LAYER M1 ;
    RECT -0.159 -0.039  0.025  0.039 ;
  LAYER V1 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V12_2x1_WEST

VIA CDS_V12_1x3_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.173  0.025  0.173 ;
  LAYER V1 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M2 ;
    RECT -0.057 -0.159  0.057  0.159 ;
END CDS_V12_1x3_CENTER

VIA CDS_V12_3x1_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.159 -0.039  0.159  0.039 ;
  LAYER V1 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M2 ;
    RECT -0.191 -0.025  0.191  0.025 ;
END CDS_V12_3x1_CENTER

VIA CDS_V12_2x2_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.096 -0.110  0.096  0.110 ;
  LAYER V1 ;
    RECT -0.096 -0.096 -0.046 -0.046 ;
    RECT -0.096  0.046 -0.046  0.096 ;
    RECT  0.046 -0.096  0.096 -0.046 ;
    RECT  0.046  0.046  0.096  0.096 ;
  LAYER M2 ;
    RECT -0.128 -0.096  0.128  0.096 ;
END CDS_V12_2x2_CENTER

VIA CDS_V12_1x2_DFM_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V1 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M2 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V12_1x2_DFM_CENTER

VIA CDS_V12_1x2_DFM_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M2 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V12_1x2_DFM_NORTH

VIA CDS_V12_1x2_DFM_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V1 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V12_1x2_DFM_SOUTH

VIA CDS_V12_2x1_DFM_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V1 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M2 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V12_2x1_DFM_CENTER

VIA CDS_V12_2x1_DFM_EAST DEFAULT
  LAYER M1 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V12_2x1_DFM_EAST

VIA CDS_V12_2x1_DFM_WEST DEFAULT
  LAYER M1 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V1 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V12_2x1_DFM_WEST

VIA CDS_V12_1x1_MIN_AREA_VCENTER DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
END CDS_V12_1x1_MIN_AREA_VCENTER

VIA CDS_V12_1x1_MIN_AREA_HCENTER DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
END CDS_V12_1x1_MIN_AREA_HCENTER

VIA CDS_V12_1x1_MIN_AREA_VEAST DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.163  0.025 ;
END CDS_V12_1x1_MIN_AREA_VEAST

VIA CDS_V12_1x1_MIN_AREA_HEAST DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.163  0.025 ;
END CDS_V12_1x1_MIN_AREA_HEAST

VIA CDS_V12_1x1_MIN_AREA_VWEST DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.163 -0.025  0.057  0.025 ;
END CDS_V12_1x1_MIN_AREA_VWEST

VIA CDS_V12_1x1_MIN_AREA_HWEST DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.163 -0.025  0.057  0.025 ;
END CDS_V12_1x1_MIN_AREA_HWEST

VIA CDS_V12_1x2_S_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.033  0.033  0.167 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V12_1x2_S_NORTH

VIA CDS_V12_1x2_S_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.167  0.033  0.033 ;
  LAYER V1 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V12_1x2_S_SOUTH

VIA CDS_V12_1x2_S_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.100  0.033  0.100 ;
  LAYER V1 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M2 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V12_1x2_S_CENTER

VIA CDS_V12_1x2_S_DFM_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.033  0.033  0.167 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M2 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V12_1x2_S_DFM_NORTH

VIA CDS_V12_1x2_S_DFM_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.167  0.033  0.033 ;
  LAYER V1 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V12_1x2_S_DFM_SOUTH

VIA CDS_V12_1x2_S_DFM_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.100  0.033  0.100 ;
  LAYER V1 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M2 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V12_1x2_S_DFM_CENTER

VIA CDS_V12_2x1_S_DFM_EAST DEFAULT
  LAYER M1 ;
    RECT -0.033 -0.033  0.167  0.033 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M2 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V12_2x1_S_DFM_EAST

VIA CDS_V12_2x1_S_DFM_WEST DEFAULT
  LAYER M1 ;
    RECT -0.167 -0.033  0.033  0.033 ;
  LAYER V1 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V12_2x1_S_DFM_WEST

VIA CDS_V12_2x1_S_DFM_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.100 -0.033  0.100  0.033 ;
  LAYER V1 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M2 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V12_2x1_S_DFM_CENTER

VIA CDS_V23_1x1_VH DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V23_1x1_VH

VIA CDS_V23_1x1_VV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V23_1x1_VV

VIA CDS_V23_1x1_HH DEFAULT
  LAYER M2 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V23_1x1_HH

VIA CDS_V23_1x1_HV DEFAULT
  LAYER M2 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V23_1x1_HV

VIA CDS_V23_1x2_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.092  0.039  0.092 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V23_1x2_CENTER

VIA CDS_V23_1x2_NORTH DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.025  0.039  0.159 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V23_1x2_NORTH

VIA CDS_V23_1x2_SOUTH DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.159  0.039  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V23_1x2_SOUTH

VIA CDS_V23_2x1_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V23_2x1_CENTER

VIA CDS_V23_2x1_EAST DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V23_2x1_EAST

VIA CDS_V23_2x1_WEST DEFAULT
  LAYER M2 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V23_2x1_WEST

VIA CDS_V23_1x3_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.159  0.039  0.159 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.191 ;
END CDS_V23_1x3_CENTER

VIA CDS_V23_3x1_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.173 -0.025  0.173  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.159 -0.057  0.159  0.057 ;
END CDS_V23_3x1_CENTER

VIA CDS_V23_2x2_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.110 -0.096  0.110  0.096 ;
  LAYER V2 ;
    RECT -0.096 -0.096 -0.046 -0.046 ;
    RECT -0.096  0.046 -0.046  0.096 ;
    RECT  0.046 -0.096  0.096 -0.046 ;
    RECT  0.046  0.046  0.096  0.096 ;
  LAYER M3 ;
    RECT -0.096 -0.128  0.096  0.128 ;
END CDS_V23_2x2_CENTER

VIA CDS_V23_1x2_DFM_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V23_1x2_DFM_CENTER

VIA CDS_V23_1x2_DFM_NORTH DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V23_1x2_DFM_NORTH

VIA CDS_V23_1x2_DFM_SOUTH DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V23_1x2_DFM_SOUTH

VIA CDS_V23_2x1_DFM_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V23_2x1_DFM_CENTER

VIA CDS_V23_2x1_DFM_EAST DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V23_2x1_DFM_EAST

VIA CDS_V23_2x1_DFM_WEST DEFAULT
  LAYER M2 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V23_2x1_DFM_WEST

VIA CDS_V23_1x1_MIN_AREA_C_V DEFAULT
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V23_1x1_MIN_AREA_C_V

VIA CDS_V23_1x1_MIN_AREA_E_V DEFAULT
  LAYER M2 ;
    RECT -0.042 -0.025  0.178  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V23_1x1_MIN_AREA_E_V

VIA CDS_V23_1x1_MIN_AREA_W_V DEFAULT
  LAYER M2 ;
    RECT -0.178 -0.025  0.042  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V23_1x1_MIN_AREA_W_V

VIA CDS_V23_2x1_MIN_AREA_E_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V23_2x1_MIN_AREA_E_EASTH

VIA CDS_V23_2x1_MIN_AREA_E_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V23_2x1_MIN_AREA_E_WESTH

VIA CDS_V23_2x1_MIN_AREA_C_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V23_2x1_MIN_AREA_C_EASTH

VIA CDS_V23_2x1_MIN_AREA_C_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V23_2x1_MIN_AREA_C_WESTH

VIA CDS_V23_2x1_MIN_AREA_W_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V23_2x1_MIN_AREA_W_EASTH

VIA CDS_V23_2x1_MIN_AREA_W_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V23_2x1_MIN_AREA_W_WESTH

VIA CDS_V23_1x2_MIN_AREA_N_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V23_1x2_MIN_AREA_N_NORTHV

VIA CDS_V23_1x2_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V23_1x2_MIN_AREA_N_SOUTHV

VIA CDS_V23_1x2_MIN_AREA_C_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V23_1x2_MIN_AREA_C_NORTHV

VIA CDS_V23_1x2_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V23_1x2_MIN_AREA_C_SOUTHV

VIA CDS_V23_1x2_MIN_AREA_S_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V23_1x2_MIN_AREA_S_NORTHV

VIA CDS_V23_1x2_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V23_1x2_MIN_AREA_S_SOUTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_N_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V23_1x2_DFM_MIN_AREA_N_NORTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V23_1x2_DFM_MIN_AREA_N_SOUTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_C_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V23_1x2_DFM_MIN_AREA_C_NORTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V23_1x2_DFM_MIN_AREA_C_SOUTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_S_NORTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M3 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V23_1x2_DFM_MIN_AREA_S_NORTHV

VIA CDS_V23_1x2_DFM_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V2 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V23_1x2_DFM_MIN_AREA_S_SOUTHV

VIA CDS_V23_2x1_DFM_MIN_AREA_E_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_E_EASTH

VIA CDS_V23_2x1_DFM_MIN_AREA_E_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_E_WESTH

VIA CDS_V23_2x1_DFM_MIN_AREA_C_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_C_EASTH

VIA CDS_V23_2x1_DFM_MIN_AREA_C_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_C_WESTH

VIA CDS_V23_2x1_DFM_MIN_AREA_W_EASTH DEFAULT
  LAYER M2 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M3 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_W_EASTH

VIA CDS_V23_2x1_DFM_MIN_AREA_W_WESTH DEFAULT
  LAYER M2 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V2 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M3 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_W_WESTH

VIA CDS_V23_1x2_MIN_AREA_C_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V23_1x2_MIN_AREA_C_VCENTER

VIA CDS_V23_1x2_MIN_AREA_N_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V23_1x2_MIN_AREA_N_VCENTER

VIA CDS_V23_1x2_MIN_AREA_S_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V23_1x2_MIN_AREA_S_VCENTER

VIA CDS_V23_1x2_DFM_MIN_AREA_C_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V23_1x2_DFM_MIN_AREA_C_VCENTER

VIA CDS_V23_1x2_DFM_MIN_AREA_N_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V23_1x2_DFM_MIN_AREA_N_VCENTER

VIA CDS_V23_1x2_DFM_MIN_AREA_S_VCENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V23_1x2_DFM_MIN_AREA_S_VCENTER

VIA CDS_V23_2x1_DFM_MIN_AREA_C_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_C_HCENTER

VIA CDS_V23_2x1_DFM_MIN_AREA_E_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_E_HCENTER

VIA CDS_V23_2x1_DFM_MIN_AREA_W_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V23_2x1_DFM_MIN_AREA_W_HCENTER

VIA CDS_V23_2x1_MIN_AREA_C_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V23_2x1_MIN_AREA_C_HCENTER

VIA CDS_V23_2x1_MIN_AREA_E_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V23_2x1_MIN_AREA_E_HCENTER

VIA CDS_V23_2x1_MIN_AREA_W_HCENTER DEFAULT
  LAYER M2 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V23_2x1_MIN_AREA_W_HCENTER

VIA CDS_V34_1x1_VH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V34_1x1_VH

VIA CDS_V34_1x1_VV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V34_1x1_VV

VIA CDS_V34_1x1_HH DEFAULT
  LAYER M3 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V34_1x1_HH

VIA CDS_V34_1x1_HV DEFAULT
  LAYER M3 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V34_1x1_HV

VIA CDS_V34_1x2_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V34_1x2_CENTER

VIA CDS_V34_1x2_NORTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V34_1x2_NORTH

VIA CDS_V34_1x2_SOUTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V34_1x2_SOUTH

VIA CDS_V34_2x1_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.092 -0.039  0.092  0.039 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V34_2x1_CENTER

VIA CDS_V34_2x1_EAST DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.039  0.159  0.039 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V34_2x1_EAST

VIA CDS_V34_2x1_WEST DEFAULT
  LAYER M3 ;
    RECT -0.159 -0.039  0.025  0.039 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V34_2x1_WEST

VIA CDS_V34_1x3_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.173  0.025  0.173 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.057 -0.159  0.057  0.159 ;
END CDS_V34_1x3_CENTER

VIA CDS_V34_3x1_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.159 -0.039  0.159  0.039 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.191  0.025 ;
END CDS_V34_3x1_CENTER

VIA CDS_V34_2x2_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.096 -0.110  0.096  0.110 ;
  LAYER V3 ;
    RECT -0.096 -0.096 -0.046 -0.046 ;
    RECT -0.096  0.046 -0.046  0.096 ;
    RECT  0.046 -0.096  0.096 -0.046 ;
    RECT  0.046  0.046  0.096  0.096 ;
  LAYER M4 ;
    RECT -0.128 -0.096  0.128  0.096 ;
END CDS_V34_2x2_CENTER

VIA CDS_V34_1x2_DFM_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V34_1x2_DFM_CENTER

VIA CDS_V34_1x2_DFM_NORTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V34_1x2_DFM_NORTH

VIA CDS_V34_1x2_DFM_SOUTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V34_1x2_DFM_SOUTH

VIA CDS_V34_2x1_DFM_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V34_2x1_DFM_CENTER

VIA CDS_V34_2x1_DFM_EAST DEFAULT
  LAYER M3 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V34_2x1_DFM_EAST

VIA CDS_V34_2x1_DFM_WEST DEFAULT
  LAYER M3 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V34_2x1_DFM_WEST

VIA CDS_V34_1x1_MIN_AREA_C_H DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V34_1x1_MIN_AREA_C_H

VIA CDS_V34_1x1_MIN_AREA_N_H DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.042  0.025  0.178 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V34_1x1_MIN_AREA_N_H

VIA CDS_V34_1x1_MIN_AREA_S_H DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.178  0.025  0.042 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V34_1x1_MIN_AREA_S_H

VIA CDS_V34_2x1_MIN_AREA_E_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V34_2x1_MIN_AREA_E_EASTH

VIA CDS_V34_2x1_MIN_AREA_E_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V34_2x1_MIN_AREA_E_WESTH

VIA CDS_V34_2x1_MIN_AREA_C_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V34_2x1_MIN_AREA_C_EASTH

VIA CDS_V34_2x1_MIN_AREA_C_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V34_2x1_MIN_AREA_C_WESTH

VIA CDS_V34_2x1_MIN_AREA_W_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V34_2x1_MIN_AREA_W_EASTH

VIA CDS_V34_2x1_MIN_AREA_W_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V34_2x1_MIN_AREA_W_WESTH

VIA CDS_V34_1x2_MIN_AREA_N_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V34_1x2_MIN_AREA_N_NORTHV

VIA CDS_V34_1x2_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V34_1x2_MIN_AREA_N_SOUTHV

VIA CDS_V34_1x2_MIN_AREA_C_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V34_1x2_MIN_AREA_C_NORTHV

VIA CDS_V34_1x2_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V34_1x2_MIN_AREA_C_SOUTHV

VIA CDS_V34_1x2_MIN_AREA_S_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V34_1x2_MIN_AREA_S_NORTHV

VIA CDS_V34_1x2_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V34_1x2_MIN_AREA_S_SOUTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_N_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V34_1x2_DFM_MIN_AREA_N_NORTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V34_1x2_DFM_MIN_AREA_N_SOUTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_C_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V34_1x2_DFM_MIN_AREA_C_NORTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V34_1x2_DFM_MIN_AREA_C_SOUTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_S_NORTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M4 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V34_1x2_DFM_MIN_AREA_S_NORTHV

VIA CDS_V34_1x2_DFM_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V3 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V34_1x2_DFM_MIN_AREA_S_SOUTHV

VIA CDS_V34_2x1_DFM_MIN_AREA_E_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_E_EASTH

VIA CDS_V34_2x1_DFM_MIN_AREA_E_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_E_WESTH

VIA CDS_V34_2x1_DFM_MIN_AREA_C_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_C_EASTH

VIA CDS_V34_2x1_DFM_MIN_AREA_C_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_C_WESTH

VIA CDS_V34_2x1_DFM_MIN_AREA_W_EASTH DEFAULT
  LAYER M3 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M4 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_W_EASTH

VIA CDS_V34_2x1_DFM_MIN_AREA_W_WESTH DEFAULT
  LAYER M3 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V3 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M4 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_W_WESTH

VIA CDS_V34_1x2_MIN_AREA_C_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V34_1x2_MIN_AREA_C_VCENTER

VIA CDS_V34_1x2_MIN_AREA_N_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V34_1x2_MIN_AREA_N_VCENTER

VIA CDS_V34_1x2_MIN_AREA_S_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V34_1x2_MIN_AREA_S_VCENTER

VIA CDS_V34_1x2_DFM_MIN_AREA_C_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V34_1x2_DFM_MIN_AREA_C_VCENTER

VIA CDS_V34_1x2_DFM_MIN_AREA_N_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V34_1x2_DFM_MIN_AREA_N_VCENTER

VIA CDS_V34_1x2_DFM_MIN_AREA_S_VCENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V34_1x2_DFM_MIN_AREA_S_VCENTER

VIA CDS_V34_2x1_DFM_MIN_AREA_C_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_C_HCENTER

VIA CDS_V34_2x1_DFM_MIN_AREA_E_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_E_HCENTER

VIA CDS_V34_2x1_DFM_MIN_AREA_W_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V34_2x1_DFM_MIN_AREA_W_HCENTER

VIA CDS_V34_2x1_MIN_AREA_C_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V34_2x1_MIN_AREA_C_HCENTER

VIA CDS_V34_2x1_MIN_AREA_E_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V34_2x1_MIN_AREA_E_HCENTER

VIA CDS_V34_2x1_MIN_AREA_W_HCENTER DEFAULT
  LAYER M3 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V34_2x1_MIN_AREA_W_HCENTER

VIA CDS_V45_1x1_VH DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V45_1x1_VH

VIA CDS_V45_1x1_VV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V45_1x1_VV

VIA CDS_V45_1x1_HH DEFAULT
  LAYER M4 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V45_1x1_HH

VIA CDS_V45_1x1_HV DEFAULT
  LAYER M4 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V45_1x1_HV

VIA CDS_V45_1x2_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.092  0.039  0.092 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V45_1x2_CENTER

VIA CDS_V45_1x2_NORTH DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.025  0.039  0.159 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V45_1x2_NORTH

VIA CDS_V45_1x2_SOUTH DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.159  0.039  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V45_1x2_SOUTH

VIA CDS_V45_2x1_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V45_2x1_CENTER

VIA CDS_V45_2x1_EAST DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V45_2x1_EAST

VIA CDS_V45_2x1_WEST DEFAULT
  LAYER M4 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V45_2x1_WEST

VIA CDS_V45_1x3_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.159  0.039  0.159 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.191 ;
END CDS_V45_1x3_CENTER

VIA CDS_V45_3x1_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.173 -0.025  0.173  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.159 -0.057  0.159  0.057 ;
END CDS_V45_3x1_CENTER

VIA CDS_V45_2x2_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.110 -0.096  0.110  0.096 ;
  LAYER V4 ;
    RECT -0.096 -0.096 -0.046 -0.046 ;
    RECT -0.096  0.046 -0.046  0.096 ;
    RECT  0.046 -0.096  0.096 -0.046 ;
    RECT  0.046  0.046  0.096  0.096 ;
  LAYER M5 ;
    RECT -0.096 -0.128  0.096  0.128 ;
END CDS_V45_2x2_CENTER

VIA CDS_V45_1x2_DFM_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V45_1x2_DFM_CENTER

VIA CDS_V45_1x2_DFM_NORTH DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V45_1x2_DFM_NORTH

VIA CDS_V45_1x2_DFM_SOUTH DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V45_1x2_DFM_SOUTH

VIA CDS_V45_2x1_DFM_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V45_2x1_DFM_CENTER

VIA CDS_V45_2x1_DFM_EAST DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V45_2x1_DFM_EAST

VIA CDS_V45_2x1_DFM_WEST DEFAULT
  LAYER M4 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V45_2x1_DFM_WEST

VIA CDS_V45_1x1_MIN_AREA_C_V DEFAULT
  LAYER M4 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V45_1x1_MIN_AREA_C_V

VIA CDS_V45_1x1_MIN_AREA_E_V DEFAULT
  LAYER M4 ;
    RECT -0.042 -0.025  0.178  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V45_1x1_MIN_AREA_E_V

VIA CDS_V45_1x1_MIN_AREA_W_V DEFAULT
  LAYER M4 ;
    RECT -0.178 -0.025  0.042  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V45_1x1_MIN_AREA_W_V

VIA CDS_V45_2x1_MIN_AREA_E_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V45_2x1_MIN_AREA_E_EASTH

VIA CDS_V45_2x1_MIN_AREA_E_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V45_2x1_MIN_AREA_E_WESTH

VIA CDS_V45_2x1_MIN_AREA_C_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V45_2x1_MIN_AREA_C_EASTH

VIA CDS_V45_2x1_MIN_AREA_C_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V45_2x1_MIN_AREA_C_WESTH

VIA CDS_V45_2x1_MIN_AREA_W_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V45_2x1_MIN_AREA_W_EASTH

VIA CDS_V45_2x1_MIN_AREA_W_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V45_2x1_MIN_AREA_W_WESTH

VIA CDS_V45_1x2_MIN_AREA_N_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V45_1x2_MIN_AREA_N_NORTHV

VIA CDS_V45_1x2_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V45_1x2_MIN_AREA_N_SOUTHV

VIA CDS_V45_1x2_MIN_AREA_C_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V45_1x2_MIN_AREA_C_NORTHV

VIA CDS_V45_1x2_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V45_1x2_MIN_AREA_C_SOUTHV

VIA CDS_V45_1x2_MIN_AREA_S_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V45_1x2_MIN_AREA_S_NORTHV

VIA CDS_V45_1x2_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V45_1x2_MIN_AREA_S_SOUTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_N_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V45_1x2_DFM_MIN_AREA_N_NORTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V45_1x2_DFM_MIN_AREA_N_SOUTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_C_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V45_1x2_DFM_MIN_AREA_C_NORTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V45_1x2_DFM_MIN_AREA_C_SOUTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_S_NORTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M5 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V45_1x2_DFM_MIN_AREA_S_NORTHV

VIA CDS_V45_1x2_DFM_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V4 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V45_1x2_DFM_MIN_AREA_S_SOUTHV

VIA CDS_V45_2x1_DFM_MIN_AREA_E_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_E_EASTH

VIA CDS_V45_2x1_DFM_MIN_AREA_E_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_E_WESTH

VIA CDS_V45_2x1_DFM_MIN_AREA_C_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_C_EASTH

VIA CDS_V45_2x1_DFM_MIN_AREA_C_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_C_WESTH

VIA CDS_V45_2x1_DFM_MIN_AREA_W_EASTH DEFAULT
  LAYER M4 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M5 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_W_EASTH

VIA CDS_V45_2x1_DFM_MIN_AREA_W_WESTH DEFAULT
  LAYER M4 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V4 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M5 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_W_WESTH

VIA CDS_V45_1x2_MIN_AREA_C_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V45_1x2_MIN_AREA_C_VCENTER

VIA CDS_V45_1x2_MIN_AREA_N_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V45_1x2_MIN_AREA_N_VCENTER

VIA CDS_V45_1x2_MIN_AREA_S_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V45_1x2_MIN_AREA_S_VCENTER

VIA CDS_V45_1x2_DFM_MIN_AREA_C_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V45_1x2_DFM_MIN_AREA_C_VCENTER

VIA CDS_V45_1x2_DFM_MIN_AREA_N_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V45_1x2_DFM_MIN_AREA_N_VCENTER

VIA CDS_V45_1x2_DFM_MIN_AREA_S_VCENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V45_1x2_DFM_MIN_AREA_S_VCENTER

VIA CDS_V45_2x1_DFM_MIN_AREA_C_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_C_HCENTER

VIA CDS_V45_2x1_DFM_MIN_AREA_E_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_E_HCENTER

VIA CDS_V45_2x1_DFM_MIN_AREA_W_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V45_2x1_DFM_MIN_AREA_W_HCENTER

VIA CDS_V45_2x1_MIN_AREA_C_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V45_2x1_MIN_AREA_C_HCENTER

VIA CDS_V45_2x1_MIN_AREA_E_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V45_2x1_MIN_AREA_E_HCENTER

VIA CDS_V45_2x1_MIN_AREA_W_HCENTER DEFAULT
  LAYER M4 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V45_2x1_MIN_AREA_W_HCENTER

VIA CDS_V56_1x1_VH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V56_1x1_VH

VIA CDS_V56_1x1_VV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.042  0.025  0.042 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V56_1x1_VV

VIA CDS_V56_1x1_HH DEFAULT
  LAYER M5 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V56_1x1_HH

VIA CDS_V56_1x1_HV DEFAULT
  LAYER M5 ;
    RECT -0.042 -0.025  0.042  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.057 ;
END CDS_V56_1x1_HV

VIA CDS_V56_1x2_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V56_1x2_CENTER

VIA CDS_V56_1x2_NORTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V56_1x2_NORTH

VIA CDS_V56_1x2_SOUTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V56_1x2_SOUTH

VIA CDS_V56_2x1_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.092 -0.039  0.092  0.039 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V56_2x1_CENTER

VIA CDS_V56_2x1_EAST DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.039  0.159  0.039 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V56_2x1_EAST

VIA CDS_V56_2x1_WEST DEFAULT
  LAYER M5 ;
    RECT -0.159 -0.039  0.025  0.039 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V56_2x1_WEST

VIA CDS_V56_1x3_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.173  0.025  0.173 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.057 -0.159  0.057  0.159 ;
END CDS_V56_1x3_CENTER

VIA CDS_V56_3x1_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.159 -0.039  0.159  0.039 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.191  0.025 ;
END CDS_V56_3x1_CENTER

VIA CDS_V56_2x2_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.096 -0.110  0.096  0.110 ;
  LAYER V5 ;
    RECT -0.096 -0.096 -0.046 -0.046 ;
    RECT -0.096  0.046 -0.046  0.096 ;
    RECT  0.046 -0.096  0.096 -0.046 ;
    RECT  0.046  0.046  0.096  0.096 ;
  LAYER M6 ;
    RECT -0.128 -0.096  0.128  0.096 ;
END CDS_V56_2x2_CENTER

VIA CDS_V56_1x2_DFM_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.106  0.025  0.106 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V56_1x2_DFM_CENTER

VIA CDS_V56_1x2_DFM_NORTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.039  0.025  0.173 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V56_1x2_DFM_NORTH

VIA CDS_V56_1x2_DFM_SOUTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.173  0.025  0.039 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V56_1x2_DFM_SOUTH

VIA CDS_V56_2x1_DFM_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.106 -0.025  0.106  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V56_2x1_DFM_CENTER

VIA CDS_V56_2x1_DFM_EAST DEFAULT
  LAYER M5 ;
    RECT -0.039 -0.025  0.173  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V56_2x1_DFM_EAST

VIA CDS_V56_2x1_DFM_WEST DEFAULT
  LAYER M5 ;
    RECT -0.173 -0.025  0.039  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V56_2x1_DFM_WEST

VIA CDS_V56_1x1_MIN_AREA_C_H DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V56_1x1_MIN_AREA_C_H

VIA CDS_V56_1x1_MIN_AREA_N_H DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.042  0.025  0.178 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V56_1x1_MIN_AREA_N_H

VIA CDS_V56_1x1_MIN_AREA_S_H DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.178  0.025  0.042 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.025 ;
END CDS_V56_1x1_MIN_AREA_S_H

VIA CDS_V56_2x1_MIN_AREA_E_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V56_2x1_MIN_AREA_E_EASTH

VIA CDS_V56_2x1_MIN_AREA_E_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V56_2x1_MIN_AREA_E_WESTH

VIA CDS_V56_2x1_MIN_AREA_C_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V56_2x1_MIN_AREA_C_EASTH

VIA CDS_V56_2x1_MIN_AREA_C_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V56_2x1_MIN_AREA_C_WESTH

VIA CDS_V56_2x1_MIN_AREA_W_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.159  0.057 ;
END CDS_V56_2x1_MIN_AREA_W_EASTH

VIA CDS_V56_2x1_MIN_AREA_W_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.159 -0.057  0.025  0.057 ;
END CDS_V56_2x1_MIN_AREA_W_WESTH

VIA CDS_V56_1x2_MIN_AREA_N_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V56_1x2_MIN_AREA_N_NORTHV

VIA CDS_V56_1x2_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V56_1x2_MIN_AREA_N_SOUTHV

VIA CDS_V56_1x2_MIN_AREA_C_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V56_1x2_MIN_AREA_C_NORTHV

VIA CDS_V56_1x2_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V56_1x2_MIN_AREA_C_SOUTHV

VIA CDS_V56_1x2_MIN_AREA_S_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.057  0.159 ;
END CDS_V56_1x2_MIN_AREA_S_NORTHV

VIA CDS_V56_1x2_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.159  0.057  0.025 ;
END CDS_V56_1x2_MIN_AREA_S_SOUTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_N_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.039  0.025  0.181 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V56_1x2_DFM_MIN_AREA_N_NORTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_N_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.173  0.025  0.047 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V56_1x2_DFM_MIN_AREA_N_SOUTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_C_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.043  0.025  0.177 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V56_1x2_DFM_MIN_AREA_C_NORTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_C_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.177  0.025  0.043 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V56_1x2_DFM_MIN_AREA_C_SOUTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_S_NORTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.047  0.025  0.173 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT -0.025  0.109  0.025  0.159 ;
  LAYER M6 ;
    RECT -0.025 -0.057  0.025  0.191 ;
END CDS_V56_1x2_DFM_MIN_AREA_S_NORTHV

VIA CDS_V56_1x2_DFM_MIN_AREA_S_SOUTHV DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.181  0.025  0.039 ;
  LAYER V5 ;
    RECT -0.025 -0.159  0.025 -0.109 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.191  0.025  0.057 ;
END CDS_V56_1x2_DFM_MIN_AREA_S_SOUTHV

VIA CDS_V56_2x1_DFM_MIN_AREA_E_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.039 -0.025  0.181  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_E_EASTH

VIA CDS_V56_2x1_DFM_MIN_AREA_E_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.173 -0.025  0.047  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_E_WESTH

VIA CDS_V56_2x1_DFM_MIN_AREA_C_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.043 -0.025  0.177  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_C_EASTH

VIA CDS_V56_2x1_DFM_MIN_AREA_C_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.177 -0.025  0.043  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_C_WESTH

VIA CDS_V56_2x1_DFM_MIN_AREA_W_EASTH DEFAULT
  LAYER M5 ;
    RECT -0.047 -0.025  0.173  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.025  0.025  0.025 ;
    RECT  0.109 -0.025  0.159  0.025 ;
  LAYER M6 ;
    RECT -0.057 -0.025  0.191  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_W_EASTH

VIA CDS_V56_2x1_DFM_MIN_AREA_W_WESTH DEFAULT
  LAYER M5 ;
    RECT -0.181 -0.025  0.039  0.025 ;
  LAYER V5 ;
    RECT -0.159 -0.025 -0.109  0.025 ;
    RECT -0.025 -0.025  0.025  0.025 ;
  LAYER M6 ;
    RECT -0.191 -0.025  0.057  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_W_WESTH

VIA CDS_V56_1x2_MIN_AREA_C_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V56_1x2_MIN_AREA_C_VCENTER

VIA CDS_V56_1x2_MIN_AREA_N_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V56_1x2_MIN_AREA_N_VCENTER

VIA CDS_V56_1x2_MIN_AREA_S_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.057 -0.092  0.057  0.092 ;
END CDS_V56_1x2_MIN_AREA_S_VCENTER

VIA CDS_V56_1x2_DFM_MIN_AREA_C_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V56_1x2_DFM_MIN_AREA_C_VCENTER

VIA CDS_V56_1x2_DFM_MIN_AREA_N_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.106  0.025  0.114 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V56_1x2_DFM_MIN_AREA_N_VCENTER

VIA CDS_V56_1x2_DFM_MIN_AREA_S_VCENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.114  0.025  0.106 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025 -0.042 ;
    RECT -0.025  0.042  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.124  0.025  0.124 ;
END CDS_V56_1x2_DFM_MIN_AREA_S_VCENTER

VIA CDS_V56_2x1_DFM_MIN_AREA_C_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_C_HCENTER

VIA CDS_V56_2x1_DFM_MIN_AREA_E_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_E_HCENTER

VIA CDS_V56_2x1_DFM_MIN_AREA_W_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.124 -0.025  0.124  0.025 ;
END CDS_V56_2x1_DFM_MIN_AREA_W_HCENTER

VIA CDS_V56_2x1_MIN_AREA_C_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V56_2x1_MIN_AREA_C_HCENTER

VIA CDS_V56_2x1_MIN_AREA_E_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.106 -0.025  0.114  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V56_2x1_MIN_AREA_E_HCENTER

VIA CDS_V56_2x1_MIN_AREA_W_HCENTER DEFAULT
  LAYER M5 ;
    RECT -0.114 -0.025  0.106  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025 -0.042  0.025 ;
    RECT  0.042 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.092 -0.057  0.092  0.057 ;
END CDS_V56_2x1_MIN_AREA_W_HCENTER

VIA CDS_V67_1x1_VH DEFAULT
  LAYER M6 ;
    RECT -0.050 -0.090  0.050  0.090 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V67_1x1_VH

VIA CDS_V67_1x1_VV DEFAULT
  LAYER M6 ;
    RECT -0.050 -0.090  0.050  0.090 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.090 ;
END CDS_V67_1x1_VV

VIA CDS_V67_1x1_HH DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.050  0.090  0.050 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V67_1x1_HH

VIA CDS_V67_1x1_HV DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.050  0.090  0.050 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.090 ;
END CDS_V67_1x1_HV

VIA CDS_V67_1x2_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.150  0.090  0.150 ;
  LAYER W0 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V67_1x2_CENTER

VIA CDS_V67_1x2_NORTH DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.050  0.090  0.250 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V67_1x2_NORTH

VIA CDS_V67_1x2_SOUTH DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.250  0.090  0.050 ;
  LAYER W0 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V67_1x2_SOUTH

VIA CDS_V67_2x1_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.190 -0.050  0.190  0.050 ;
  LAYER W0 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B1 ;
    RECT -0.150 -0.090  0.150  0.090 ;
END CDS_V67_2x1_CENTER

VIA CDS_V67_2x1_EAST DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.050  0.290  0.050 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B1 ;
    RECT -0.050 -0.090  0.250  0.090 ;
END CDS_V67_2x1_EAST

VIA CDS_V67_2x1_WEST DEFAULT
  LAYER M6 ;
    RECT -0.290 -0.050  0.090  0.050 ;
  LAYER W0 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.250 -0.090  0.050  0.090 ;
END CDS_V67_2x1_WEST

VIA CDS_V67_1x3_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.250  0.090  0.250 ;
  LAYER W0 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.290 ;
END CDS_V67_1x3_CENTER

VIA CDS_V67_3x1_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.290 -0.050  0.290  0.050 ;
  LAYER W0 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B1 ;
    RECT -0.250 -0.090  0.250  0.090 ;
END CDS_V67_3x1_CENTER

VIA CDS_V67_2x2_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.190 -0.150  0.190  0.150 ;
  LAYER W0 ;
    RECT -0.150 -0.150 -0.050 -0.050 ;
    RECT -0.150  0.050 -0.050  0.150 ;
    RECT  0.050 -0.150  0.150 -0.050 ;
    RECT  0.050  0.050  0.150  0.150 ;
  LAYER B1 ;
    RECT -0.150 -0.190  0.150  0.190 ;
END CDS_V67_2x2_CENTER

VIA CDS_V67_1x2_DFM_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.050 -0.190  0.050  0.190 ;
  LAYER W0 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V67_1x2_DFM_CENTER

VIA CDS_V67_1x2_DFM_NORTH DEFAULT
  LAYER M6 ;
    RECT -0.050 -0.090  0.050  0.290 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V67_1x2_DFM_NORTH

VIA CDS_V67_1x2_DFM_SOUTH DEFAULT
  LAYER M6 ;
    RECT -0.050 -0.290  0.050  0.090 ;
  LAYER W0 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V67_1x2_DFM_SOUTH

VIA CDS_V67_2x1_DFM_CENTER DEFAULT
  LAYER M6 ;
    RECT -0.190 -0.050  0.190  0.050 ;
  LAYER W0 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B1 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V67_2x1_DFM_CENTER

VIA CDS_V67_2x1_DFM_EAST DEFAULT
  LAYER M6 ;
    RECT -0.090 -0.050  0.290  0.050 ;
  LAYER W0 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B1 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V67_2x1_DFM_EAST

VIA CDS_V67_2x1_DFM_WEST DEFAULT
  LAYER M6 ;
    RECT -0.290 -0.050  0.090  0.050 ;
  LAYER W0 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B1 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V67_2x1_DFM_WEST

VIA CDS_V78_1x1_VH DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V78_1x1_VH

VIA CDS_V78_1x1_VV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.090 ;
END CDS_V78_1x1_VV

VIA CDS_V78_1x1_HH DEFAULT
  LAYER B1 ;
    RECT -0.090 -0.050  0.090  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V78_1x1_HH

VIA CDS_V78_1x1_HV DEFAULT
  LAYER B1 ;
    RECT -0.090 -0.050  0.090  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.090 ;
END CDS_V78_1x1_HV

VIA CDS_V78_1x2_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.190 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.090 -0.150  0.090  0.150 ;
END CDS_V78_1x2_CENTER

VIA CDS_V78_1x2_NORTH DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.290 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.250 ;
END CDS_V78_1x2_NORTH

VIA CDS_V78_1x2_SOUTH DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.250  0.090  0.050 ;
END CDS_V78_1x2_SOUTH

VIA CDS_V78_2x1_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.150 -0.090  0.150  0.090 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V78_2x1_CENTER

VIA CDS_V78_2x1_EAST DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.250  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V78_2x1_EAST

VIA CDS_V78_2x1_WEST DEFAULT
  LAYER B1 ;
    RECT -0.250 -0.090  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V78_2x1_WEST

VIA CDS_V78_1x3_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.290 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.090 -0.250  0.090  0.250 ;
END CDS_V78_1x3_CENTER

VIA CDS_V78_3x1_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.250 -0.090  0.250  0.090 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.290  0.050 ;
END CDS_V78_3x1_CENTER

VIA CDS_V78_2x2_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.150 -0.190  0.150  0.190 ;
  LAYER W1 ;
    RECT -0.150 -0.150 -0.050 -0.050 ;
    RECT -0.150  0.050 -0.050  0.150 ;
    RECT  0.050 -0.150  0.150 -0.050 ;
    RECT  0.050  0.050  0.150  0.150 ;
  LAYER B2 ;
    RECT -0.190 -0.150  0.190  0.150 ;
END CDS_V78_2x2_CENTER

VIA CDS_V78_1x2_DFM_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.190 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V78_1x2_DFM_CENTER

VIA CDS_V78_1x2_DFM_NORTH DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.290 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V78_1x2_DFM_NORTH

VIA CDS_V78_1x2_DFM_SOUTH DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V78_1x2_DFM_SOUTH

VIA CDS_V78_2x1_DFM_CENTER DEFAULT
  LAYER B1 ;
    RECT -0.190 -0.050  0.190  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V78_2x1_DFM_CENTER

VIA CDS_V78_2x1_DFM_EAST DEFAULT
  LAYER B1 ;
    RECT -0.090 -0.050  0.290  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V78_2x1_DFM_EAST

VIA CDS_V78_2x1_DFM_WEST DEFAULT
  LAYER B1 ;
    RECT -0.290 -0.050  0.090  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V78_2x1_DFM_WEST

VIA CDS_V78_1x1_MIN_AREA_C_H DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.200  0.050  0.200 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V78_1x1_MIN_AREA_C_H

VIA CDS_V78_1x1_MIN_AREA_N_H DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.310 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V78_1x1_MIN_AREA_N_H

VIA CDS_V78_1x1_MIN_AREA_S_H DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.310  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.050 ;
END CDS_V78_1x1_MIN_AREA_S_H

VIA CDS_V78_2x1_MIN_AREA_E_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.090 -0.050  0.310  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.250  0.090 ;
END CDS_V78_2x1_MIN_AREA_E_EASTH

VIA CDS_V78_2x1_MIN_AREA_E_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.290 -0.050  0.110  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.250 -0.090  0.050  0.090 ;
END CDS_V78_2x1_MIN_AREA_E_WESTH

VIA CDS_V78_2x1_MIN_AREA_C_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.100 -0.050  0.300  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.250  0.090 ;
END CDS_V78_2x1_MIN_AREA_C_EASTH

VIA CDS_V78_2x1_MIN_AREA_C_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.300 -0.050  0.100  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.250 -0.090  0.050  0.090 ;
END CDS_V78_2x1_MIN_AREA_C_WESTH

VIA CDS_V78_2x1_MIN_AREA_W_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.110 -0.050  0.290  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.250  0.090 ;
END CDS_V78_2x1_MIN_AREA_W_EASTH

VIA CDS_V78_2x1_MIN_AREA_W_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.310 -0.050  0.090  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.250 -0.090  0.050  0.090 ;
END CDS_V78_2x1_MIN_AREA_W_WESTH

VIA CDS_V78_1x2_MIN_AREA_N_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.310 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.250 ;
END CDS_V78_1x2_MIN_AREA_N_NORTHV

VIA CDS_V78_1x2_MIN_AREA_N_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.110 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.250  0.090  0.050 ;
END CDS_V78_1x2_MIN_AREA_N_SOUTHV

VIA CDS_V78_1x2_MIN_AREA_C_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.100  0.050  0.300 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.250 ;
END CDS_V78_1x2_MIN_AREA_C_NORTHV

VIA CDS_V78_1x2_MIN_AREA_C_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.300  0.050  0.100 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.250  0.090  0.050 ;
END CDS_V78_1x2_MIN_AREA_C_SOUTHV

VIA CDS_V78_1x2_MIN_AREA_S_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.110  0.050  0.290 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.090  0.250 ;
END CDS_V78_1x2_MIN_AREA_S_NORTHV

VIA CDS_V78_1x2_MIN_AREA_S_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.310  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.250  0.090  0.050 ;
END CDS_V78_1x2_MIN_AREA_S_SOUTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_N_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.090  0.050  0.310 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V78_1x2_DFM_MIN_AREA_N_NORTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_N_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.290  0.050  0.110 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V78_1x2_DFM_MIN_AREA_N_SOUTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_C_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.100  0.050  0.300 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V78_1x2_DFM_MIN_AREA_C_NORTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_C_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.300  0.050  0.100 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V78_1x2_DFM_MIN_AREA_C_SOUTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_S_NORTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.110  0.050  0.290 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT -0.050  0.150  0.050  0.250 ;
  LAYER B2 ;
    RECT -0.050 -0.090  0.050  0.290 ;
END CDS_V78_1x2_DFM_MIN_AREA_S_NORTHV

VIA CDS_V78_1x2_DFM_MIN_AREA_S_SOUTHV DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.310  0.050  0.090 ;
  LAYER W1 ;
    RECT -0.050 -0.250  0.050 -0.150 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.050 -0.290  0.050  0.090 ;
END CDS_V78_1x2_DFM_MIN_AREA_S_SOUTHV

VIA CDS_V78_2x1_DFM_MIN_AREA_E_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.090 -0.050  0.310  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_E_EASTH

VIA CDS_V78_2x1_DFM_MIN_AREA_E_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.290 -0.050  0.110  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_E_WESTH

VIA CDS_V78_2x1_DFM_MIN_AREA_C_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.100 -0.050  0.300  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_C_EASTH

VIA CDS_V78_2x1_DFM_MIN_AREA_C_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.300 -0.050  0.100  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_C_WESTH

VIA CDS_V78_2x1_DFM_MIN_AREA_W_EASTH DEFAULT
  LAYER B1 ;
    RECT -0.110 -0.050  0.290  0.050 ;
  LAYER W1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
    RECT  0.150 -0.050  0.250  0.050 ;
  LAYER B2 ;
    RECT -0.090 -0.050  0.290  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_W_EASTH

VIA CDS_V78_2x1_DFM_MIN_AREA_W_WESTH DEFAULT
  LAYER B1 ;
    RECT -0.310 -0.050  0.090  0.050 ;
  LAYER W1 ;
    RECT -0.250 -0.050 -0.150  0.050 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER B2 ;
    RECT -0.290 -0.050  0.090  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_W_WESTH

VIA CDS_V78_1x2_MIN_AREA_C_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.200  0.050  0.200 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.090 -0.150  0.090  0.150 ;
END CDS_V78_1x2_MIN_AREA_C_VCENTER

VIA CDS_V78_1x2_MIN_AREA_N_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.210 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.090 -0.150  0.090  0.150 ;
END CDS_V78_1x2_MIN_AREA_N_VCENTER

VIA CDS_V78_1x2_MIN_AREA_S_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.210  0.050  0.190 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.090 -0.150  0.090  0.150 ;
END CDS_V78_1x2_MIN_AREA_S_VCENTER

VIA CDS_V78_1x2_DFM_MIN_AREA_C_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.200  0.050  0.200 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V78_1x2_DFM_MIN_AREA_C_VCENTER

VIA CDS_V78_1x2_DFM_MIN_AREA_N_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.190  0.050  0.210 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V78_1x2_DFM_MIN_AREA_N_VCENTER

VIA CDS_V78_1x2_DFM_MIN_AREA_S_VCENTER DEFAULT
  LAYER B1 ;
    RECT -0.050 -0.210  0.050  0.190 ;
  LAYER W1 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT -0.050  0.050  0.050  0.150 ;
  LAYER B2 ;
    RECT -0.050 -0.190  0.050  0.190 ;
END CDS_V78_1x2_DFM_MIN_AREA_S_VCENTER

VIA CDS_V78_2x1_DFM_MIN_AREA_C_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.200 -0.050  0.200  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_C_HCENTER

VIA CDS_V78_2x1_DFM_MIN_AREA_E_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.190 -0.050  0.210  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_E_HCENTER

VIA CDS_V78_2x1_DFM_MIN_AREA_W_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.210 -0.050  0.190  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.190 -0.050  0.190  0.050 ;
END CDS_V78_2x1_DFM_MIN_AREA_W_HCENTER

VIA CDS_V78_2x1_MIN_AREA_C_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.200 -0.050  0.200  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.150 -0.090  0.150  0.090 ;
END CDS_V78_2x1_MIN_AREA_C_HCENTER

VIA CDS_V78_2x1_MIN_AREA_E_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.190 -0.050  0.210  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.150 -0.090  0.150  0.090 ;
END CDS_V78_2x1_MIN_AREA_E_HCENTER

VIA CDS_V78_2x1_MIN_AREA_W_HCENTER DEFAULT
  LAYER B1 ;
    RECT -0.210 -0.050  0.190  0.050 ;
  LAYER W1 ;
    RECT -0.150 -0.050 -0.050  0.050 ;
    RECT  0.050 -0.050  0.150  0.050 ;
  LAYER B2 ;
    RECT -0.150 -0.090  0.150  0.090 ;
END CDS_V78_2x1_MIN_AREA_W_HCENTER

VIA CDS_V89_1x1_VH DEFAULT
  LAYER B2 ;
    RECT -0.200 -0.260  0.200  0.260 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.260 -0.200  0.260  0.200 ;
END CDS_V89_1x1_VH

VIA CDS_V89_1x1_VV DEFAULT
  LAYER B2 ;
    RECT -0.200 -0.260  0.200  0.260 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.200 -0.260  0.200  0.260 ;
END CDS_V89_1x1_VV

VIA CDS_V89_1x1_HH DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.200  0.260  0.200 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.260 -0.200  0.260  0.200 ;
END CDS_V89_1x1_HH

VIA CDS_V89_1x1_HV DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.200  0.260  0.200 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.200 -0.260  0.200  0.260 ;
END CDS_V89_1x1_HV

VIA CDS_V89_1x2_CENTER DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.600  0.260  0.600 ;
  LAYER YZ ;
    RECT -0.180 -0.580  0.180 -0.220 ;
    RECT -0.180  0.220  0.180  0.580 ;
  LAYER IA ;
    RECT -0.200 -0.660  0.200  0.660 ;
END CDS_V89_1x2_CENTER

VIA CDS_V89_1x2_NORTH DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.200  0.260  1.000 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT -0.180  0.620  0.180  0.980 ;
  LAYER IA ;
    RECT -0.200 -0.260  0.200  1.060 ;
END CDS_V89_1x2_NORTH

VIA CDS_V89_1x2_SOUTH DEFAULT
  LAYER B2 ;
    RECT -0.260 -1.000  0.260  0.200 ;
  LAYER YZ ;
    RECT -0.180 -0.980  0.180 -0.620 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.200 -1.060  0.200  0.260 ;
END CDS_V89_1x2_SOUTH

VIA CDS_V89_2x1_CENTER DEFAULT
  LAYER B2 ;
    RECT -0.660 -0.200  0.660  0.200 ;
  LAYER YZ ;
    RECT -0.580 -0.180 -0.220  0.180 ;
    RECT  0.220 -0.180  0.580  0.180 ;
  LAYER IA ;
    RECT -0.600 -0.260  0.600  0.260 ;
END CDS_V89_2x1_CENTER

VIA CDS_V89_2x1_EAST DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.200  1.060  0.200 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT  0.620 -0.180  0.980  0.180 ;
  LAYER IA ;
    RECT -0.200 -0.260  1.000  0.260 ;
END CDS_V89_2x1_EAST

VIA CDS_V89_2x1_WEST DEFAULT
  LAYER B2 ;
    RECT -1.060 -0.200  0.260  0.200 ;
  LAYER YZ ;
    RECT -0.980 -0.180 -0.620  0.180 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -1.000 -0.260  0.200  0.260 ;
END CDS_V89_2x1_WEST

VIA CDS_V89_1x2_DFM_CENTER DEFAULT
  LAYER B2 ;
    RECT -0.200 -0.660  0.200  0.660 ;
  LAYER YZ ;
    RECT -0.180 -0.580  0.180 -0.220 ;
    RECT -0.180  0.220  0.180  0.580 ;
  LAYER IA ;
    RECT -0.200 -0.660  0.200  0.660 ;
END CDS_V89_1x2_DFM_CENTER

VIA CDS_V89_1x2_DFM_NORTH DEFAULT
  LAYER B2 ;
    RECT -0.200 -0.260  0.200  1.060 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT -0.180  0.620  0.180  0.980 ;
  LAYER IA ;
    RECT -0.200 -0.260  0.200  1.060 ;
END CDS_V89_1x2_DFM_NORTH

VIA CDS_V89_1x2_DFM_SOUTH DEFAULT
  LAYER B2 ;
    RECT -0.200 -1.060  0.200  0.260 ;
  LAYER YZ ;
    RECT -0.180 -0.980  0.180 -0.620 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -0.200 -1.060  0.200  0.260 ;
END CDS_V89_1x2_DFM_SOUTH

VIA CDS_V89_2x1_DFM_CENTER DEFAULT
  LAYER B2 ;
    RECT -0.660 -0.200  0.660  0.200 ;
  LAYER YZ ;
    RECT -0.580 -0.180 -0.220  0.180 ;
    RECT  0.220 -0.180  0.580  0.180 ;
  LAYER IA ;
    RECT -0.660 -0.200  0.660  0.200 ;
END CDS_V89_2x1_DFM_CENTER

VIA CDS_V89_2x1_DFM_EAST DEFAULT
  LAYER B2 ;
    RECT -0.260 -0.200  1.060  0.200 ;
  LAYER YZ ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT  0.620 -0.180  0.980  0.180 ;
  LAYER IA ;
    RECT -0.260 -0.200  1.060  0.200 ;
END CDS_V89_2x1_DFM_EAST

VIA CDS_V89_2x1_DFM_WEST DEFAULT
  LAYER B2 ;
    RECT -1.060 -0.200  0.260  0.200 ;
  LAYER YZ ;
    RECT -0.980 -0.180 -0.620  0.180 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IA ;
    RECT -1.060 -0.200  0.260  0.200 ;
END CDS_V89_2x1_DFM_WEST

VIA CDS_V910_1x1_VH DEFAULT
  LAYER IA ;
    RECT -0.200 -0.260  0.200  0.260 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -0.260 -0.200  0.260  0.200 ;
END CDS_V910_1x1_VH

VIA CDS_V910_1x1_VV DEFAULT
  LAYER IA ;
    RECT -0.200 -0.260  0.200  0.260 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -0.200 -0.260  0.200  0.260 ;
END CDS_V910_1x1_VV

VIA CDS_V910_1x1_HH DEFAULT
  LAYER IA ;
    RECT -0.260 -0.200  0.260  0.200 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -0.260 -0.200  0.260  0.200 ;
END CDS_V910_1x1_HH

VIA CDS_V910_1x1_HV DEFAULT
  LAYER IA ;
    RECT -0.260 -0.200  0.260  0.200 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -0.200 -0.260  0.200  0.260 ;
END CDS_V910_1x1_HV

VIA CDS_V910_1x2_CENTER DEFAULT
  LAYER IA ;
    RECT -0.260 -0.600  0.260  0.600 ;
  LAYER XA ;
    RECT -0.180 -0.580  0.180 -0.220 ;
    RECT -0.180  0.220  0.180  0.580 ;
  LAYER IB ;
    RECT -0.200 -0.660  0.200  0.660 ;
END CDS_V910_1x2_CENTER

VIA CDS_V910_1x2_NORTH DEFAULT
  LAYER IA ;
    RECT -0.260 -0.200  0.260  1.000 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT -0.180  0.620  0.180  0.980 ;
  LAYER IB ;
    RECT -0.200 -0.260  0.200  1.060 ;
END CDS_V910_1x2_NORTH

VIA CDS_V910_1x2_SOUTH DEFAULT
  LAYER IA ;
    RECT -0.260 -1.000  0.260  0.200 ;
  LAYER XA ;
    RECT -0.180 -0.980  0.180 -0.620 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -0.200 -1.060  0.200  0.260 ;
END CDS_V910_1x2_SOUTH

VIA CDS_V910_2x1_CENTER DEFAULT
  LAYER IA ;
    RECT -0.660 -0.200  0.660  0.200 ;
  LAYER XA ;
    RECT -0.580 -0.180 -0.220  0.180 ;
    RECT  0.220 -0.180  0.580  0.180 ;
  LAYER IB ;
    RECT -0.600 -0.260  0.600  0.260 ;
END CDS_V910_2x1_CENTER

VIA CDS_V910_2x1_EAST DEFAULT
  LAYER IA ;
    RECT -0.260 -0.200  1.060  0.200 ;
  LAYER XA ;
    RECT -0.180 -0.180  0.180  0.180 ;
    RECT  0.620 -0.180  0.980  0.180 ;
  LAYER IB ;
    RECT -0.200 -0.260  1.000  0.260 ;
END CDS_V910_2x1_EAST

VIA CDS_V910_2x1_WEST DEFAULT
  LAYER IA ;
    RECT -1.060 -0.200  0.260  0.200 ;
  LAYER XA ;
    RECT -0.980 -0.180 -0.620  0.180 ;
    RECT -0.180 -0.180  0.180  0.180 ;
  LAYER IB ;
    RECT -1.000 -0.260  0.200  0.260 ;
END CDS_V910_2x1_WEST

VIA CDS_V1011_1x1_VH DEFAULT
  LAYER IB ;
    RECT -2.000 -2.000  2.000  2.000 ;
  LAYER VV ;
    RECT -1.500 -1.500  1.500  1.500 ;
  LAYER LB ;
    RECT -2.500 -2.500  2.500  2.500 ;
END CDS_V1011_1x1_VH

################################ END VIA FOR ROUTING ####################################

################################ VIA BAR FOR ROUTING ####################################

# "Standard" VxBAR

VIA CDS_V12_BAR_H_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V1 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M2 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V12_BAR_H_CENTER

VIA CDS_V12_BAR_H_EAST DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.092  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.075  0.025 ;
  LAYER M2 ;
    RECT -0.042 -0.025  0.092  0.025 ;
END CDS_V12_BAR_H_EAST

VIA CDS_V12_BAR_H_WEST DEFAULT
  LAYER M1 ;
    RECT -0.092 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.075 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.092 -0.025  0.042  0.025 ;
END CDS_V12_BAR_H_WEST

VIA CDS_V12_BAR_V_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.067  0.025  0.067 ;
  LAYER V1 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M2 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V12_BAR_V_CENTER

VIA CDS_V12_BAR_V_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.042  0.025  0.092 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.025  0.075 ;
  LAYER M2 ;
    RECT -0.025 -0.042  0.025  0.092 ;
END CDS_V12_BAR_V_NORTH

VIA CDS_V12_BAR_V_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.092  0.025  0.042 ;
  LAYER V1 ;
    RECT -0.025 -0.075  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.092  0.025  0.042 ;
END CDS_V12_BAR_V_SOUTH

VIA CDS_V23_BAR_H_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V2 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M3 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V23_BAR_H_CENTER

VIA CDS_V23_BAR_V_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.067  0.025  0.067 ;
  LAYER V2 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M3 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V23_BAR_V_CENTER

VIA CDS_V34_BAR_H_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V3 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M4 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V34_BAR_H_CENTER

VIA CDS_V34_BAR_V_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.067  0.025  0.067 ;
  LAYER V3 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M4 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V34_BAR_V_CENTER

VIA CDS_V45_BAR_H_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V4 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M5 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V45_BAR_H_CENTER

VIA CDS_V45_BAR_V_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.067  0.025  0.067 ;
  LAYER V4 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M5 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V45_BAR_V_CENTER

VIA CDS_V56_BAR_H_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V5 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M6 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V56_BAR_H_CENTER

VIA CDS_V56_BAR_V_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.067  0.025  0.067 ;
  LAYER V5 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M6 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V56_BAR_V_CENTER

# "Shifted" VxBAR

VIA CDS_V12_BAR_SHIFTED_H_EAST DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V1 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V12_BAR_SHIFTED_H_EAST

VIA CDS_V12_BAR_SHIFTED_H_WEST DEFAULT
  LAYER M1 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V1 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M2 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V12_BAR_SHIFTED_H_WEST

VIA CDS_V12_BAR_SHIFTED_V_NORTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.025  0.025  0.109 ;
  LAYER V1 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M2 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V12_BAR_SHIFTED_V_NORTH

VIA CDS_V12_BAR_SHIFTED_V_SOUTH DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.109  0.025  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M2 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V12_BAR_SHIFTED_V_SOUTH

VIA CDS_V23_BAR_SHIFTED_H_EAST DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V2 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V23_BAR_SHIFTED_H_EAST

VIA CDS_V23_BAR_SHIFTED_H_WEST DEFAULT
  LAYER M2 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M3 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V23_BAR_SHIFTED_H_WEST

VIA CDS_V23_BAR_SHIFTED_V_NORTH DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.025  0.025  0.109 ;
  LAYER V2 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M3 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V23_BAR_SHIFTED_V_NORTH

VIA CDS_V23_BAR_SHIFTED_V_SOUTH DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.109  0.025  0.025 ;
  LAYER V2 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M3 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V23_BAR_SHIFTED_V_SOUTH

VIA CDS_V34_BAR_SHIFTED_H_EAST DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V3 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M4 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V34_BAR_SHIFTED_H_EAST

VIA CDS_V34_BAR_SHIFTED_H_WEST DEFAULT
  LAYER M3 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V3 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M4 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V34_BAR_SHIFTED_H_WEST

VIA CDS_V34_BAR_SHIFTED_V_NORTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.025  0.025  0.109 ;
  LAYER V3 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V34_BAR_SHIFTED_V_NORTH

VIA CDS_V34_BAR_SHIFTED_V_SOUTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.109  0.025  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M4 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V34_BAR_SHIFTED_V_SOUTH

VIA CDS_V45_BAR_SHIFTED_H_EAST DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V4 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V45_BAR_SHIFTED_H_EAST

VIA CDS_V45_BAR_SHIFTED_H_WEST DEFAULT
  LAYER M4 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M5 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V45_BAR_SHIFTED_H_WEST

VIA CDS_V45_BAR_SHIFTED_V_NORTH DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.025  0.025  0.109 ;
  LAYER V4 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M5 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V45_BAR_SHIFTED_V_NORTH

VIA CDS_V45_BAR_SHIFTED_V_SOUTH DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.109  0.025  0.025 ;
  LAYER V4 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M5 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V45_BAR_SHIFTED_V_SOUTH

VIA CDS_V56_BAR_SHIFTED_H_EAST DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V5 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M6 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V56_BAR_SHIFTED_H_EAST

VIA CDS_V56_BAR_SHIFTED_H_WEST DEFAULT
  LAYER M5 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V5 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M6 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V56_BAR_SHIFTED_H_WEST

VIA CDS_V56_BAR_SHIFTED_V_NORTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.025  0.025  0.109 ;
  LAYER V5 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V56_BAR_SHIFTED_V_NORTH

VIA CDS_V56_BAR_SHIFTED_V_SOUTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.109  0.025  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M6 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V56_BAR_SHIFTED_V_SOUTH

# "Standard min area" VxBAR
#    V12: top layer only
#    V23 and above: bottom layer only

VIA CDS_V12_BAR_MIN_AREA_H_CENTER DEFAULT
  LAYER M1 ;
    RECT -0.067 -0.025  0.067  0.025 ;
  LAYER V1 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
END CDS_V12_BAR_MIN_AREA_H_CENTER

VIA CDS_V12_BAR_MIN_AREA_H_EAST DEFAULT
  LAYER M1 ;
    RECT -0.042 -0.025  0.092  0.025 ;
  LAYER V1 ;
    RECT -0.025 -0.025  0.075  0.025 ;
  LAYER M2 ;
    RECT -0.042 -0.025  0.178  0.025 ;
END CDS_V12_BAR_MIN_AREA_H_EAST

VIA CDS_V12_BAR_MIN_AREA_H_WEST DEFAULT
  LAYER M1 ;
    RECT -0.092 -0.025  0.042  0.025 ;
  LAYER V1 ;
    RECT -0.075 -0.025  0.025  0.025 ;
  LAYER M2 ;
    RECT -0.178 -0.025  0.042  0.025 ;
END CDS_V12_BAR_MIN_AREA_H_WEST

VIA CDS_V23_BAR_MIN_AREA_H_CENTER DEFAULT
  LAYER M2 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V2 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M3 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V23_BAR_MIN_AREA_H_CENTER

VIA CDS_V34_BAR_MIN_AREA_V_CENTER DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V3 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M4 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V34_BAR_MIN_AREA_V_CENTER

VIA CDS_V45_BAR_MIN_AREA_H_CENTER DEFAULT
  LAYER M4 ;
    RECT -0.110 -0.025  0.110  0.025 ;
  LAYER V4 ;
    RECT -0.050 -0.025  0.050  0.025 ;
  LAYER M5 ;
    RECT -0.067 -0.025  0.067  0.025 ;
END CDS_V45_BAR_MIN_AREA_H_CENTER

VIA CDS_V56_BAR_MIN_AREA_V_CENTER DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.110  0.025  0.110 ;
  LAYER V5 ;
    RECT -0.025 -0.050  0.025  0.050 ;
  LAYER M6 ;
    RECT -0.025 -0.067  0.025  0.067 ;
END CDS_V56_BAR_MIN_AREA_V_CENTER

# "Shifted min area" VxBAR
#    V12: top layer only
#    V23 and above: bottom layer only

VIA CDS_V12_BAR_MIN_AREA_SHIFTED_H_EAST DEFAULT
  LAYER M1 ;
    RECT -0.025 -0.025  0.109  0.025 ;
  LAYER V1 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.025  0.195  0.025 ;
END CDS_V12_BAR_MIN_AREA_SHIFTED_H_EAST

VIA CDS_V12_BAR_MIN_AREA_SHIFTED_H_WEST DEFAULT
  LAYER M1 ;
    RECT -0.109 -0.025  0.025  0.025 ;
  LAYER V1 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M2 ;
    RECT -0.195 -0.025  0.025  0.025 ;
END CDS_V12_BAR_MIN_AREA_SHIFTED_H_WEST

VIA CDS_V23_BAR_MIN_AREA_SHIFTED_H_EAST DEFAULT
  LAYER M2 ;
    RECT -0.025 -0.025  0.195  0.025 ;
  LAYER V2 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V23_BAR_MIN_AREA_SHIFTED_H_EAST

VIA CDS_V23_BAR_MIN_AREA_SHIFTED_H_WEST DEFAULT
  LAYER M2 ;
    RECT -0.195 -0.025  0.025  0.025 ;
  LAYER V2 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M3 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V23_BAR_MIN_AREA_SHIFTED_H_WEST

VIA CDS_V34_BAR_MIN_AREA_SHIFTED_V_NORTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.025  0.025  0.195 ;
  LAYER V3 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M4 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V34_BAR_MIN_AREA_SHIFTED_V_NORTH

VIA CDS_V34_BAR_MIN_AREA_SHIFTED_V_SOUTH DEFAULT
  LAYER M3 ;
    RECT -0.025 -0.195  0.025  0.025 ;
  LAYER V3 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M4 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V34_BAR_MIN_AREA_SHIFTED_V_SOUTH

VIA CDS_V45_BAR_MIN_AREA_SHIFTED_H_EAST DEFAULT
  LAYER M4 ;
    RECT -0.025 -0.025  0.195  0.025 ;
  LAYER V4 ;
    RECT -0.008 -0.025  0.092  0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.025  0.109  0.025 ;
END CDS_V45_BAR_MIN_AREA_SHIFTED_H_EAST

VIA CDS_V45_BAR_MIN_AREA_SHIFTED_H_WEST DEFAULT
  LAYER M4 ;
    RECT -0.195 -0.025  0.025  0.025 ;
  LAYER V4 ;
    RECT -0.092 -0.025  0.008  0.025 ;
  LAYER M5 ;
    RECT -0.109 -0.025  0.025  0.025 ;
END CDS_V45_BAR_MIN_AREA_SHIFTED_H_WEST

VIA CDS_V56_BAR_MIN_AREA_SHIFTED_V_NORTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.025  0.025  0.195 ;
  LAYER V5 ;
    RECT -0.025 -0.008  0.025  0.092 ;
  LAYER M6 ;
    RECT -0.025 -0.025  0.025  0.109 ;
END CDS_V56_BAR_MIN_AREA_SHIFTED_V_NORTH

VIA CDS_V56_BAR_MIN_AREA_SHIFTED_V_SOUTH DEFAULT
  LAYER M5 ;
    RECT -0.025 -0.195  0.025  0.025 ;
  LAYER V5 ;
    RECT -0.025 -0.092  0.025  0.008 ;
  LAYER M6 ;
    RECT -0.025 -0.109  0.025  0.025 ;
END CDS_V56_BAR_MIN_AREA_SHIFTED_V_SOUTH

############################## END VIA BAR FOR ROUTING ##################################

################################ VIA LRG FOR ROUTING ####################################

VIA CDS_V12_LRG
  LAYER M1 ;
    RECT -0.067 -0.067  0.067  0.067 ;
  LAYER V1 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER M2 ;
    RECT -0.082 -0.082  0.082  0.082 ;
END CDS_V12_LRG

VIA CDS_V23_LRG
  LAYER M2 ;
    RECT -0.082 -0.082  0.082  0.082 ;
  LAYER V2 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER M3 ;
    RECT -0.082 -0.082  0.082  0.082 ;
END CDS_V23_LRG

VIA CDS_V34_LRG
  LAYER M3 ;
    RECT -0.082 -0.082  0.082  0.082 ;
  LAYER V3 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER M4 ;
    RECT -0.082 -0.082  0.082  0.082 ;
END CDS_V34_LRG

VIA CDS_V45_LRG
  LAYER M4 ;
    RECT -0.082 -0.082  0.082  0.082 ;
  LAYER V4 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER M5 ;
    RECT -0.082 -0.082  0.082  0.082 ;
END CDS_V45_LRG

VIA CDS_V56_LRG
  LAYER M5 ;
    RECT -0.082 -0.082  0.082  0.082 ;
  LAYER V5 ;
    RECT -0.050 -0.050  0.050  0.050 ;
  LAYER M6 ;
    RECT -0.082 -0.082  0.082  0.082 ;
END CDS_V56_LRG

############################## END VIA LRG FOR ROUTING ##################################

END LIBRARY
